magic
tech sky130A
magscale 1 2
timestamp 1698166509
<< obsli1 >>
rect 1104 2159 138828 137649
<< obsm1 >>
rect 14 2128 138828 137680
<< metal2 >>
rect 5142 139200 5254 139800
rect 10938 139200 11050 139800
rect 16734 139200 16846 139800
rect 23174 139200 23286 139800
rect 28970 139200 29082 139800
rect 34766 139200 34878 139800
rect 41206 139200 41318 139800
rect 47002 139200 47114 139800
rect 52798 139200 52910 139800
rect 59238 139200 59350 139800
rect 65034 139200 65146 139800
rect 70830 139200 70942 139800
rect 77270 139200 77382 139800
rect 83066 139200 83178 139800
rect 88862 139200 88974 139800
rect 95302 139200 95414 139800
rect 101098 139200 101210 139800
rect 106894 139200 107006 139800
rect 113334 139200 113446 139800
rect 119130 139200 119242 139800
rect 124926 139200 125038 139800
rect 131366 139200 131478 139800
rect 137162 139200 137274 139800
rect -10 200 102 800
rect 5786 200 5898 800
rect 11582 200 11694 800
rect 17378 200 17490 800
rect 23818 200 23930 800
rect 29614 200 29726 800
rect 35410 200 35522 800
rect 41850 200 41962 800
rect 47646 200 47758 800
rect 53442 200 53554 800
rect 59882 200 59994 800
rect 65678 200 65790 800
rect 71474 200 71586 800
rect 77914 200 78026 800
rect 83710 200 83822 800
rect 89506 200 89618 800
rect 95946 200 96058 800
rect 101742 200 101854 800
rect 107538 200 107650 800
rect 113978 200 114090 800
rect 119774 200 119886 800
rect 125570 200 125682 800
rect 132010 200 132122 800
rect 137806 200 137918 800
<< obsm2 >>
rect 20 139856 138626 139890
rect 20 139144 5086 139856
rect 5310 139144 10882 139856
rect 11106 139144 16678 139856
rect 16902 139144 23118 139856
rect 23342 139144 28914 139856
rect 29138 139144 34710 139856
rect 34934 139144 41150 139856
rect 41374 139144 46946 139856
rect 47170 139144 52742 139856
rect 52966 139144 59182 139856
rect 59406 139144 64978 139856
rect 65202 139144 70774 139856
rect 70998 139144 77214 139856
rect 77438 139144 83010 139856
rect 83234 139144 88806 139856
rect 89030 139144 95246 139856
rect 95470 139144 101042 139856
rect 101266 139144 106838 139856
rect 107062 139144 113278 139856
rect 113502 139144 119074 139856
rect 119298 139144 124870 139856
rect 125094 139144 131310 139856
rect 131534 139144 137106 139856
rect 137330 139144 138626 139856
rect 20 856 138626 139144
rect 158 800 5730 856
rect 5954 800 11526 856
rect 11750 800 17322 856
rect 17546 800 23762 856
rect 23986 800 29558 856
rect 29782 800 35354 856
rect 35578 800 41794 856
rect 42018 800 47590 856
rect 47814 800 53386 856
rect 53610 800 59826 856
rect 60050 800 65622 856
rect 65846 800 71418 856
rect 71642 800 77858 856
rect 78082 800 83654 856
rect 83878 800 89450 856
rect 89674 800 95890 856
rect 96114 800 101686 856
rect 101910 800 107482 856
rect 107706 800 113922 856
rect 114146 800 119718 856
rect 119942 800 125514 856
rect 125738 800 131954 856
rect 132178 800 137750 856
rect 137974 800 138626 856
<< metal3 >>
rect 200 139348 800 139588
rect 139200 136628 139800 136914
rect 200 132548 800 132788
rect 139200 130508 139800 130748
rect 200 126428 800 126668
rect 139200 123662 139800 123948
rect 200 120308 800 120548
rect 139200 117542 139800 117828
rect 200 113508 800 113748
rect 139200 111468 139800 111754
rect 200 107388 800 107628
rect 139200 104622 139800 104908
rect 200 101268 800 101508
rect 139200 98548 139800 98834
rect 200 94468 800 94708
rect 139200 92428 139800 92714
rect 200 88348 800 88588
rect 139200 85582 139800 85868
rect 200 82228 800 82468
rect 139200 79508 139800 79794
rect 200 75428 800 75668
rect 139200 73388 139800 73674
rect 200 69308 800 69548
rect 139200 66588 139800 66874
rect 200 63188 800 63428
rect 139200 60422 139800 60708
rect 200 56388 800 56628
rect 139200 54348 139800 54588
rect 200 50268 800 50508
rect 139200 47502 139800 47788
rect 200 44148 800 44388
rect 139200 41382 139800 41668
rect 200 37348 800 37588
rect 139200 35308 139800 35594
rect 200 31228 800 31468
rect 139200 28508 139800 28794
rect 200 25108 800 25348
rect 139200 22388 139800 22674
rect 200 18308 800 18548
rect 139200 16268 139800 16508
rect 200 12188 800 12428
rect 139200 9422 139800 9708
rect 200 6068 800 6308
rect 139200 3348 139800 3588
<< obsm3 >>
rect 880 139268 139962 139501
rect 800 136994 139962 139268
rect 800 136548 139120 136994
rect 139880 136548 139962 136994
rect 800 132868 139962 136548
rect 880 132468 139962 132868
rect 800 130828 139962 132468
rect 800 130428 139120 130828
rect 139880 130428 139962 130828
rect 800 126748 139962 130428
rect 880 126348 139962 126748
rect 800 124028 139962 126348
rect 800 123582 139120 124028
rect 139880 123582 139962 124028
rect 800 120628 139962 123582
rect 880 120228 139962 120628
rect 800 117908 139962 120228
rect 800 117462 139120 117908
rect 139880 117462 139962 117908
rect 800 113828 139962 117462
rect 880 113428 139962 113828
rect 800 111834 139962 113428
rect 800 111388 139120 111834
rect 139880 111388 139962 111834
rect 800 107708 139962 111388
rect 880 107308 139962 107708
rect 800 104988 139962 107308
rect 800 104542 139120 104988
rect 139880 104542 139962 104988
rect 800 101588 139962 104542
rect 880 101188 139962 101588
rect 800 98914 139962 101188
rect 800 98468 139120 98914
rect 139880 98468 139962 98914
rect 800 94788 139962 98468
rect 880 94388 139962 94788
rect 800 92794 139962 94388
rect 800 92348 139120 92794
rect 139880 92348 139962 92794
rect 800 88668 139962 92348
rect 880 88268 139962 88668
rect 800 85948 139962 88268
rect 800 85502 139120 85948
rect 139880 85502 139962 85948
rect 800 82548 139962 85502
rect 880 82148 139962 82548
rect 800 79874 139962 82148
rect 800 79428 139120 79874
rect 139880 79428 139962 79874
rect 800 75748 139962 79428
rect 880 75348 139962 75748
rect 800 73754 139962 75348
rect 800 73308 139120 73754
rect 139880 73308 139962 73754
rect 800 69628 139962 73308
rect 880 69228 139962 69628
rect 800 66954 139962 69228
rect 800 66508 139120 66954
rect 139880 66508 139962 66954
rect 800 63508 139962 66508
rect 880 63108 139962 63508
rect 800 60788 139962 63108
rect 800 60342 139120 60788
rect 139880 60342 139962 60788
rect 800 56708 139962 60342
rect 880 56308 139962 56708
rect 800 54668 139962 56308
rect 800 54268 139120 54668
rect 139880 54268 139962 54668
rect 800 50588 139962 54268
rect 880 50188 139962 50588
rect 800 47868 139962 50188
rect 800 47422 139120 47868
rect 139880 47422 139962 47868
rect 800 44468 139962 47422
rect 880 44068 139962 44468
rect 800 41748 139962 44068
rect 800 41302 139120 41748
rect 139880 41302 139962 41748
rect 800 37668 139962 41302
rect 880 37268 139962 37668
rect 800 35674 139962 37268
rect 800 35228 139120 35674
rect 139880 35228 139962 35674
rect 800 31548 139962 35228
rect 880 31148 139962 31548
rect 800 28874 139962 31148
rect 800 28428 139120 28874
rect 139880 28428 139962 28874
rect 800 25428 139962 28428
rect 880 25028 139962 25428
rect 800 22754 139962 25028
rect 800 22308 139120 22754
rect 139880 22308 139962 22754
rect 800 18628 139962 22308
rect 880 18228 139962 18628
rect 800 16588 139962 18228
rect 800 16188 139120 16588
rect 139880 16188 139962 16588
rect 800 12508 139962 16188
rect 880 12108 139962 12508
rect 800 9788 139962 12108
rect 800 9342 139120 9788
rect 139880 9342 139962 9788
rect 800 6388 139962 9342
rect 880 5988 139962 6388
rect 800 3668 139962 5988
rect 800 3268 139120 3668
rect 139880 3268 139962 3668
rect 800 2143 139962 3268
<< metal4 >>
rect 4208 2128 4528 137680
rect 19568 2128 19888 137680
rect 34928 2128 35248 137680
rect 50288 2128 50608 137680
rect 65648 2128 65968 137680
rect 81008 2128 81328 137680
rect 96368 2128 96688 137680
rect 111728 2128 112048 137680
rect 127088 2128 127408 137680
<< obsm4 >>
rect 31523 2347 34848 137325
rect 35328 2347 50208 137325
rect 50688 2347 65568 137325
rect 66048 2347 80928 137325
rect 81408 2347 96288 137325
rect 96768 2347 111261 137325
<< labels >>
rlabel metal3 s 200 12188 800 12428 6 i_clk
port 1 nsew signal input
rlabel metal2 s 131366 139200 131478 139800 6 i_debug_map_overlay
port 2 nsew signal input
rlabel metal3 s 200 63188 800 63428 6 i_debug_trace_overlay
port 3 nsew signal input
rlabel metal2 s 125570 200 125682 800 6 i_debug_vec_overlay
port 4 nsew signal input
rlabel metal2 s 52798 139200 52910 139800 6 i_gpout0_sel[0]
port 5 nsew signal input
rlabel metal2 s 59238 139200 59350 139800 6 i_gpout0_sel[1]
port 6 nsew signal input
rlabel metal2 s 65034 139200 65146 139800 6 i_gpout0_sel[2]
port 7 nsew signal input
rlabel metal2 s 53442 200 53554 800 6 i_gpout0_sel[3]
port 8 nsew signal input
rlabel metal3 s 139200 28508 139800 28794 6 i_gpout0_sel[4]
port 9 nsew signal input
rlabel metal2 s 124926 139200 125038 139800 6 i_gpout0_sel[5]
port 10 nsew signal input
rlabel metal2 s 77270 139200 77382 139800 6 i_gpout1_sel[0]
port 11 nsew signal input
rlabel metal2 s 47646 200 47758 800 6 i_gpout1_sel[1]
port 12 nsew signal input
rlabel metal3 s 139200 41382 139800 41668 6 i_gpout1_sel[2]
port 13 nsew signal input
rlabel metal3 s 139200 60422 139800 60708 6 i_gpout1_sel[3]
port 14 nsew signal input
rlabel metal3 s 139200 123662 139800 123948 6 i_gpout1_sel[4]
port 15 nsew signal input
rlabel metal3 s 139200 111468 139800 111754 6 i_gpout1_sel[5]
port 16 nsew signal input
rlabel metal3 s 139200 16268 139800 16508 6 i_gpout2_sel[0]
port 17 nsew signal input
rlabel metal3 s 200 101268 800 101508 6 i_gpout2_sel[1]
port 18 nsew signal input
rlabel metal2 s 29614 200 29726 800 6 i_gpout2_sel[2]
port 19 nsew signal input
rlabel metal3 s 139200 92428 139800 92714 6 i_gpout2_sel[3]
port 20 nsew signal input
rlabel metal3 s 200 107388 800 107628 6 i_gpout2_sel[4]
port 21 nsew signal input
rlabel metal3 s 200 50268 800 50508 6 i_gpout2_sel[5]
port 22 nsew signal input
rlabel metal3 s 139200 98548 139800 98834 6 i_gpout3_sel[0]
port 23 nsew signal input
rlabel metal2 s 132010 200 132122 800 6 i_gpout3_sel[1]
port 24 nsew signal input
rlabel metal2 s 88862 139200 88974 139800 6 i_gpout3_sel[2]
port 25 nsew signal input
rlabel metal2 s 5142 139200 5254 139800 6 i_gpout3_sel[3]
port 26 nsew signal input
rlabel metal3 s 139200 104622 139800 104908 6 i_gpout3_sel[4]
port 27 nsew signal input
rlabel metal3 s 200 69308 800 69548 6 i_gpout3_sel[5]
port 28 nsew signal input
rlabel metal3 s 200 82228 800 82468 6 i_gpout4_sel[0]
port 29 nsew signal input
rlabel metal3 s 200 6068 800 6308 6 i_gpout4_sel[1]
port 30 nsew signal input
rlabel metal2 s 107538 200 107650 800 6 i_gpout4_sel[2]
port 31 nsew signal input
rlabel metal3 s 200 120308 800 120548 6 i_gpout4_sel[3]
port 32 nsew signal input
rlabel metal2 s 95302 139200 95414 139800 6 i_gpout4_sel[4]
port 33 nsew signal input
rlabel metal2 s 101098 139200 101210 139800 6 i_gpout4_sel[5]
port 34 nsew signal input
rlabel metal2 s 119774 200 119886 800 6 i_gpout5_sel[0]
port 35 nsew signal input
rlabel metal2 s 70830 139200 70942 139800 6 i_gpout5_sel[1]
port 36 nsew signal input
rlabel metal3 s 139200 117542 139800 117828 6 i_gpout5_sel[2]
port 37 nsew signal input
rlabel metal2 s 83710 200 83822 800 6 i_gpout5_sel[3]
port 38 nsew signal input
rlabel metal3 s 200 75428 800 75668 6 i_gpout5_sel[4]
port 39 nsew signal input
rlabel metal3 s 139200 3348 139800 3588 6 i_gpout5_sel[5]
port 40 nsew signal input
rlabel metal3 s 139200 54348 139800 54588 6 i_mode[0]
port 41 nsew signal input
rlabel metal3 s 200 139348 800 139588 6 i_mode[1]
port 42 nsew signal input
rlabel metal3 s 200 37348 800 37588 6 i_mode[2]
port 43 nsew signal input
rlabel metal3 s 200 113508 800 113748 6 i_reg_csb
port 44 nsew signal input
rlabel metal3 s 200 25108 800 25348 6 i_reg_mosi
port 45 nsew signal input
rlabel metal3 s 139200 130508 139800 130748 6 i_reg_sclk
port 46 nsew signal input
rlabel metal2 s 28970 139200 29082 139800 6 i_reset_lock_a
port 47 nsew signal input
rlabel metal2 s 11582 200 11694 800 6 i_reset_lock_b
port 48 nsew signal input
rlabel metal2 s 35410 200 35522 800 6 i_tex_in[0]
port 49 nsew signal input
rlabel metal2 s 113978 200 114090 800 6 i_tex_in[1]
port 50 nsew signal input
rlabel metal3 s 139200 47502 139800 47788 6 i_tex_in[2]
port 51 nsew signal input
rlabel metal3 s 139200 22388 139800 22674 6 i_tex_in[3]
port 52 nsew signal input
rlabel metal2 s 89506 200 89618 800 6 i_vec_csb
port 53 nsew signal input
rlabel metal3 s 200 132548 800 132788 6 i_vec_mosi
port 54 nsew signal input
rlabel metal2 s 137806 200 137918 800 6 i_vec_sclk
port 55 nsew signal input
rlabel metal3 s 200 31228 800 31468 6 o_gpout[0]
port 56 nsew signal output
rlabel metal3 s 139200 35308 139800 35594 6 o_gpout[1]
port 57 nsew signal output
rlabel metal3 s 200 88348 800 88588 6 o_gpout[2]
port 58 nsew signal output
rlabel metal2 s 101742 200 101854 800 6 o_gpout[3]
port 59 nsew signal output
rlabel metal3 s 139200 85582 139800 85868 6 o_gpout[4]
port 60 nsew signal output
rlabel metal2 s 41206 139200 41318 139800 6 o_gpout[5]
port 61 nsew signal output
rlabel metal2 s 23174 139200 23286 139800 6 o_hsync
port 62 nsew signal output
rlabel metal2 s 65678 200 65790 800 6 o_rgb[0]
port 63 nsew signal output
rlabel metal2 s -10 200 102 800 6 o_rgb[10]
port 64 nsew signal output
rlabel metal2 s 77914 200 78026 800 6 o_rgb[11]
port 65 nsew signal output
rlabel metal2 s 47002 139200 47114 139800 6 o_rgb[12]
port 66 nsew signal output
rlabel metal2 s 83066 139200 83178 139800 6 o_rgb[13]
port 67 nsew signal output
rlabel metal2 s 119130 139200 119242 139800 6 o_rgb[14]
port 68 nsew signal output
rlabel metal3 s 200 94468 800 94708 6 o_rgb[15]
port 69 nsew signal output
rlabel metal2 s 17378 200 17490 800 6 o_rgb[16]
port 70 nsew signal output
rlabel metal2 s 5786 200 5898 800 6 o_rgb[17]
port 71 nsew signal output
rlabel metal2 s 137162 139200 137274 139800 6 o_rgb[18]
port 72 nsew signal output
rlabel metal2 s 106894 139200 107006 139800 6 o_rgb[19]
port 73 nsew signal output
rlabel metal2 s 59882 200 59994 800 6 o_rgb[1]
port 74 nsew signal output
rlabel metal3 s 139200 136628 139800 136914 6 o_rgb[20]
port 75 nsew signal output
rlabel metal3 s 139200 9422 139800 9708 6 o_rgb[21]
port 76 nsew signal output
rlabel metal2 s 16734 139200 16846 139800 6 o_rgb[22]
port 77 nsew signal output
rlabel metal3 s 139200 73388 139800 73674 6 o_rgb[23]
port 78 nsew signal output
rlabel metal2 s 23818 200 23930 800 6 o_rgb[2]
port 79 nsew signal output
rlabel metal2 s 41850 200 41962 800 6 o_rgb[3]
port 80 nsew signal output
rlabel metal3 s 200 56388 800 56628 6 o_rgb[4]
port 81 nsew signal output
rlabel metal3 s 139200 79508 139800 79794 6 o_rgb[5]
port 82 nsew signal output
rlabel metal2 s 71474 200 71586 800 6 o_rgb[6]
port 83 nsew signal output
rlabel metal3 s 200 18308 800 18548 6 o_rgb[7]
port 84 nsew signal output
rlabel metal2 s 113334 139200 113446 139800 6 o_rgb[8]
port 85 nsew signal output
rlabel metal2 s 10938 139200 11050 139800 6 o_rgb[9]
port 86 nsew signal output
rlabel metal2 s 34766 139200 34878 139800 6 o_tex_csb
port 87 nsew signal output
rlabel metal2 s 95946 200 96058 800 6 o_tex_oeb0
port 88 nsew signal output
rlabel metal3 s 200 44148 800 44388 6 o_tex_out0
port 89 nsew signal output
rlabel metal3 s 200 126428 800 126668 6 o_tex_sclk
port 90 nsew signal output
rlabel metal3 s 139200 66588 139800 66874 6 o_vsync
port 91 nsew signal output
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 92 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 92 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 92 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 92 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 137680 6 vccd1
port 92 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 93 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 93 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 93 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 137680 6 vssd1
port 93 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 140000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 33538416
string GDS_FILE /openlane/designs/raybox-zero/runs/RUN_2023.10.24_16.49.15/results/signoff/top_ew_algofoogle.magic.gds
string GDS_START 1344532
<< end >>

