* NGSPICE file created from top_ew_algofoogle.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

.subckt top_ew_algofoogle i_clk i_debug_map_overlay i_debug_trace_overlay i_debug_vec_overlay
+ i_gpout0_sel[0] i_gpout0_sel[1] i_gpout0_sel[2] i_gpout0_sel[3] i_gpout0_sel[4]
+ i_gpout0_sel[5] i_gpout1_sel[0] i_gpout1_sel[1] i_gpout1_sel[2] i_gpout1_sel[3]
+ i_gpout1_sel[4] i_gpout1_sel[5] i_gpout2_sel[0] i_gpout2_sel[1] i_gpout2_sel[2]
+ i_gpout2_sel[3] i_gpout2_sel[4] i_gpout2_sel[5] i_gpout3_sel[0] i_gpout3_sel[1]
+ i_gpout3_sel[2] i_gpout3_sel[3] i_gpout3_sel[4] i_gpout3_sel[5] i_gpout4_sel[0]
+ i_gpout4_sel[1] i_gpout4_sel[2] i_gpout4_sel[3] i_gpout4_sel[4] i_gpout4_sel[5]
+ i_gpout5_sel[0] i_gpout5_sel[1] i_gpout5_sel[2] i_gpout5_sel[3] i_gpout5_sel[4]
+ i_gpout5_sel[5] i_mode[0] i_mode[1] i_mode[2] i_reg_csb i_reg_mosi i_reg_sclk i_reset_lock_a
+ i_reset_lock_b i_tex_in[0] i_tex_in[1] i_tex_in[2] i_tex_in[3] i_vec_csb i_vec_mosi
+ i_vec_sclk o_gpout[0] o_gpout[1] o_gpout[2] o_gpout[3] o_gpout[4] o_gpout[5] o_hsync
+ o_rgb[0] o_rgb[10] o_rgb[11] o_rgb[12] o_rgb[13] o_rgb[14] o_rgb[15] o_rgb[16] o_rgb[17]
+ o_rgb[18] o_rgb[19] o_rgb[1] o_rgb[20] o_rgb[21] o_rgb[22] o_rgb[23] o_rgb[2] o_rgb[3]
+ o_rgb[4] o_rgb[5] o_rgb[6] o_rgb[7] o_rgb[8] o_rgb[9] o_tex_csb o_tex_oeb0 o_tex_out0
+ o_tex_sclk o_vsync vccd1 vssd1
XFILLER_246_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18869_ rbzero.spi_registers.spi_counter\[3\] _02579_ _02583_ vssd1 vssd1 vccd1 vccd1
+ _02584_ sky130_fd_sc_hd__o21a_1
XFILLER_95_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20900_ net60 _00916_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20831_ _00049_ _00847_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20762_ net106 _00778_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20693_ net70 _00709_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[73\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21314_ _00337_ _01330_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21245_ _00294_ _01261_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21176_ _00225_ _01192_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20127_ _03153_ _03155_ _03154_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__o21bai_1
XFILLER_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20058_ _03128_ vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__clkinv_2
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ net9 vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__clkbuf_2
XFILLER_73_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12880_ _05405_ _05406_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__nor2b_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11831_ rbzero.tex_b1\[39\] rbzero.tex_b1\[38\] _04544_ vssd1 vssd1 vccd1 vccd1 _04545_
+ sky130_fd_sc_hd__mux2_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ rbzero.wall_tracer.stepDistY\[5\] _07221_ _07193_ vssd1 vssd1 vccd1 vccd1
+ _07222_ sky130_fd_sc_hd__mux2_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11762_ rbzero.tex_b0\[34\] _03936_ _03929_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a21o_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13501_ _06184_ _06189_ vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10713_ _03578_ vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14481_ rbzero.wall_tracer.stepDistY\[-8\] _07165_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _07166_ sky130_fd_sc_hd__mux2_1
XFILLER_159_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _03954_ _04383_ _04391_ _04408_ _04026_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__a311o_1
X_16220_ _08828_ _08830_ vssd1 vssd1 vccd1 vccd1 _08832_ sky130_fd_sc_hd__and2_1
XFILLER_224_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13432_ _06098_ _06114_ _06120_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__or3_1
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10644_ _03542_ vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16151_ _08754_ _08762_ vssd1 vssd1 vccd1 vccd1 _08763_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13363_ _06048_ _06047_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__and2b_1
XFILLER_139_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10575_ rbzero.tex_r0\[10\] rbzero.tex_r0\[9\] _03501_ vssd1 vssd1 vccd1 vccd1 _03506_
+ sky130_fd_sc_hd__mux2_1
X_15102_ _07677_ _07679_ vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12314_ _04994_ rbzero.wall_tracer.trackDistX\[11\] vssd1 vssd1 vccd1 vccd1 _05008_
+ sky130_fd_sc_hd__and2_1
XFILLER_182_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16082_ _08555_ _08556_ _08694_ vssd1 vssd1 vccd1 vccd1 _08695_ sky130_fd_sc_hd__o21a_1
XFILLER_155_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13294_ _05634_ _05982_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__nor2_1
XFILLER_142_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15033_ _07455_ _07641_ _07646_ vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__a21oi_1
X_19910_ _03113_ vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__clkinv_2
X_12245_ _04938_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__buf_6
XFILLER_194_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12176_ _04873_ net36 _04877_ _04879_ _04881_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a32o_1
X_19841_ _03107_ vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__clkinv_2
XFILLER_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11127_ _03842_ _03845_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__nor2_1
X_16984_ _09523_ _09524_ vssd1 vssd1 vccd1 vccd1 _09525_ sky130_fd_sc_hd__nor2_1
XFILLER_228_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19772_ _03784_ _03781_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__nand2_1
XFILLER_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15935_ _07900_ _08530_ _08547_ vssd1 vssd1 vccd1 vccd1 _08549_ sky130_fd_sc_hd__nand3_1
X_11058_ _03781_ _03782_ _03784_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__o21ai_1
XFILLER_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18723_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.debug_overlay.vplaneY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__nand2_1
XTAP_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18654_ _02287_ _02383_ _02384_ _02385_ vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__a31o_1
XFILLER_236_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15866_ _07471_ _08478_ _07837_ _07697_ vssd1 vssd1 vccd1 vccd1 _08480_ sky130_fd_sc_hd__a2bb2o_1
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17605_ _10038_ _10141_ vssd1 vssd1 vccd1 vccd1 _10142_ sky130_fd_sc_hd__xor2_2
X_14817_ rbzero.debug_overlay.playerX\[-8\] vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__inv_2
XFILLER_236_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18585_ _02304_ _02320_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__nor2_1
X_15797_ _08383_ _08386_ _08410_ vssd1 vssd1 vccd1 vccd1 _08411_ sky130_fd_sc_hd__nor3_1
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17536_ _07472_ _07618_ vssd1 vssd1 vccd1 vccd1 _10073_ sky130_fd_sc_hd__nor2_1
Xtop_ew_algofoogle_142 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_142/HI o_rgb[0] sky130_fd_sc_hd__conb_1
XFILLER_33_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtop_ew_algofoogle_153 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_153/HI o_rgb[13]
+ sky130_fd_sc_hd__conb_1
X_14748_ _05113_ _07360_ _07361_ _07351_ vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__o211a_1
XFILLER_127_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17467_ _09950_ _10004_ vssd1 vssd1 vccd1 vccd1 _10005_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14679_ _07313_ vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16418_ _07567_ _07712_ vssd1 vssd1 vccd1 vccd1 _09028_ sky130_fd_sc_hd__nor2_1
XFILLER_177_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19206_ rbzero.spi_registers.spi_done _02589_ _02576_ _02587_ vssd1 vssd1 vccd1 vccd1
+ _02783_ sky130_fd_sc_hd__and4b_1
XFILLER_207_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17398_ _07472_ _07618_ _08732_ _09571_ vssd1 vssd1 vccd1 vccd1 _09936_ sky130_fd_sc_hd__or4_1
XFILLER_193_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19137_ rbzero.spi_registers.got_new_vinf vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__inv_2
X_16349_ rbzero.debug_overlay.playerY\[-3\] vssd1 vssd1 vccd1 vccd1 _08960_ sky130_fd_sc_hd__clkinv_2
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19068_ _02696_ vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18019_ _01798_ _01800_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__xor2_1
XFILLER_86_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21030_ net110 _01046_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout105 net108 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__buf_2
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout116 net122 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__buf_2
XFILLER_47_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout127 net128 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout138 net139 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_2
XFILLER_234_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20814_ _00032_ _00830_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_230_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20745_ net103 _00761_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20676_ net68 _00692_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10360_ _03391_ vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10291_ _03354_ vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__clkbuf_1
X_12030_ _04078_ _03781_ _04106_ _04104_ _04717_ _04731_ vssd1 vssd1 vccd1 vccd1 _04739_
+ sky130_fd_sc_hd__mux4_1
X_21228_ _00277_ _01244_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21159_ _00208_ _01175_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13981_ _05651_ _06321_ _06669_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__nand3_1
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15720_ _08298_ _08294_ _08297_ vssd1 vssd1 vccd1 vccd1 _08334_ sky130_fd_sc_hd__a21o_1
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12932_ _05604_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__clkbuf_4
XFILLER_111_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15651_ _08264_ _08262_ vssd1 vssd1 vccd1 vccd1 _08265_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12863_ _05499_ _05498_ _05549_ _05538_ _05551_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__o221a_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ rbzero.wall_tracer.visualWallDist\[-9\] _07253_ _07262_ _07263_ _07257_ vssd1
+ vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__o221a_1
XFILLER_15_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18370_ _02125_ _02126_ _02127_ vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__a21oi_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ rbzero.tex_b1\[61\] rbzero.tex_b1\[60\] _04032_ vssd1 vssd1 vccd1 vccd1 _04528_
+ sky130_fd_sc_hd__mux2_1
X_15582_ _08174_ _08195_ vssd1 vssd1 vccd1 vccd1 _08196_ sky130_fd_sc_hd__xor2_2
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _05353_ _05343_ _05346_ _05350_ _05444_ _05463_ vssd1 vssd1 vccd1 vccd1 _05483_
+ sky130_fd_sc_hd__mux4_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _09733_ _09735_ _09858_ vssd1 vssd1 vccd1 vccd1 _09860_ sky130_fd_sc_hd__a21o_1
XFILLER_15_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _07028_ _07076_ _07098_ _07133_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__a31oi_4
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ rbzero.tex_b0\[55\] _04143_ _04145_ _03930_ vssd1 vssd1 vccd1 vccd1 _04460_
+ sky130_fd_sc_hd__a31o_1
XFILLER_202_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17252_ _09698_ _09716_ _09790_ vssd1 vssd1 vccd1 vccd1 _09791_ sky130_fd_sc_hd__a21bo_1
XFILLER_175_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14464_ _07107_ _07149_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__or2_1
X_11676_ rbzero.tex_g1\[3\] _03964_ _03965_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__and3_1
XFILLER_128_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16203_ _08656_ _08657_ vssd1 vssd1 vccd1 vccd1 _08815_ sky130_fd_sc_hd__nor2_1
XFILLER_186_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13415_ _06028_ _05738_ _06102_ _06103_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__nand4_1
X_17183_ _09720_ _09721_ _09722_ _09593_ vssd1 vssd1 vccd1 vccd1 _09723_ sky130_fd_sc_hd__o22a_1
X_10627_ _03533_ vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__clkbuf_1
X_14395_ _07071_ vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__inv_2
XFILLER_139_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16134_ _08713_ _08745_ vssd1 vssd1 vccd1 vccd1 _08746_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13346_ _06032_ _06033_ _06034_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__and3_1
XFILLER_128_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10558_ rbzero.tex_r0\[18\] rbzero.tex_r0\[17\] _03490_ vssd1 vssd1 vccd1 vccd1 _03497_
+ sky130_fd_sc_hd__mux2_1
XFILLER_196_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16065_ _08676_ _08675_ vssd1 vssd1 vccd1 vccd1 _08678_ sky130_fd_sc_hd__and2b_1
XFILLER_185_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13277_ _05715_ _05638_ _05963_ _05964_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__o211ai_1
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10489_ rbzero.tex_r0\[51\] rbzero.tex_r0\[50\] _03457_ vssd1 vssd1 vccd1 vccd1 _03461_
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15016_ _07628_ _07629_ vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__and2_1
XFILLER_155_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12228_ o_vsync rbzero.wall_tracer.state\[5\] _04920_ vssd1 vssd1 vccd1 vccd1 _04926_
+ sky130_fd_sc_hd__and3_1
XFILLER_68_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19824_ _03105_ vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__clkinv_2
XFILLER_229_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12159_ net2 _04848_ _04849_ _04702_ _04865_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__a221o_1
XFILLER_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19755_ rbzero.pov.ready_buffer\[5\] _03067_ _03068_ rbzero.debug_overlay.vplaneY\[-4\]
+ _03015_ vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__a221o_1
X_16967_ rbzero.wall_tracer.trackDistX\[0\] rbzero.wall_tracer.stepDistX\[0\] vssd1
+ vssd1 vccd1 vccd1 _09509_ sky130_fd_sc_hd__or2_1
XFILLER_81_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18706_ _02427_ _02431_ _02432_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__a21oi_1
X_15918_ _07625_ _08531_ vssd1 vssd1 vccd1 vccd1 _08532_ sky130_fd_sc_hd__nor2_1
X_16898_ _09169_ _09173_ _09439_ vssd1 vssd1 vccd1 vccd1 _09440_ sky130_fd_sc_hd__a21boi_1
X_19686_ rbzero.debug_overlay.playerY\[3\] _03039_ vssd1 vssd1 vccd1 vccd1 _03043_
+ sky130_fd_sc_hd__or2_1
XFILLER_80_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15849_ _07672_ _07673_ _07379_ vssd1 vssd1 vccd1 vccd1 _08463_ sky130_fd_sc_hd__a21oi_1
X_18637_ rbzero.map_rom.i_col\[4\] _02369_ _09274_ vssd1 vssd1 vccd1 vccd1 _02370_
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18568_ _02293_ _02296_ _02294_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a21boi_1
XFILLER_224_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17519_ _07704_ _07707_ vssd1 vssd1 vccd1 vccd1 _10056_ sky130_fd_sc_hd__and2_2
X_18499_ _02218_ _02231_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__nand2_1
XFILLER_240_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20530_ net120 _00546_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_220_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20461_ net94 _00014_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20392_ net138 _00423_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_161_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21013_ net80 _01029_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_5907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11530_ rbzero.debug_overlay.facingX\[0\] _04243_ _04244_ rbzero.debug_overlay.facingX\[-1\]
+ _04247_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__a221o_1
XFILLER_169_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20728_ net100 _00744_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11461_ rbzero.tex_r1\[11\] _04142_ _04144_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__and3_1
X_20659_ net60 _00675_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13200_ _05615_ _05887_ _05888_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__and3_1
X_10412_ _03418_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__clkbuf_1
X_14180_ _06816_ _06822_ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__xor2_1
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11392_ _04110_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__clkinv_2
XFILLER_125_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13131_ _05488_ _05700_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__nand2_1
XFILLER_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10343_ rbzero.tex_r1\[53\] rbzero.tex_r1\[54\] _03377_ vssd1 vssd1 vccd1 vccd1 _03382_
+ sky130_fd_sc_hd__mux2_1
XFILLER_174_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13062_ _05747_ _05750_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__xor2_1
XFILLER_139_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10274_ rbzero.tex_b1\[22\] rbzero.tex_b1\[23\] _03344_ vssd1 vssd1 vccd1 vccd1 _03346_
+ sky130_fd_sc_hd__mux2_1
XFILLER_117_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12013_ _04717_ _04447_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__nand2_1
XFILLER_26_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17870_ _09429_ _08851_ _01529_ vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__or3b_1
XFILLER_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16821_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.stepDistX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _09364_ sky130_fd_sc_hd__nand2_1
XFILLER_120_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16752_ _05121_ vssd1 vssd1 vccd1 vccd1 _09303_ sky130_fd_sc_hd__buf_4
X_19540_ rbzero.pov.spi_buffer\[65\] rbzero.pov.spi_buffer\[66\] _02932_ vssd1 vssd1
+ vccd1 vccd1 _02939_ sky130_fd_sc_hd__mux2_1
X_13964_ _06596_ _06649_ _06652_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__a21o_1
XFILLER_24_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15703_ _08244_ _08270_ _08316_ vssd1 vssd1 vccd1 vccd1 _08317_ sky130_fd_sc_hd__a21oi_2
XFILLER_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12915_ _05538_ _05592_ _05596_ _05603_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__a31o_2
X_16683_ rbzero.traced_texa\[-12\] _09262_ _09258_ rbzero.wall_tracer.visualWallDist\[-12\]
+ vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19471_ rbzero.pov.spi_buffer\[32\] rbzero.pov.spi_buffer\[33\] _02899_ vssd1 vssd1
+ vccd1 vccd1 _02903_ sky130_fd_sc_hd__mux2_1
X_13895_ _06538_ _06546_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__and2_1
XFILLER_111_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15634_ _08193_ _08209_ vssd1 vssd1 vccd1 vccd1 _08248_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18422_ _02172_ _02173_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__or2b_1
XFILLER_179_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12846_ _05470_ _05447_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__nor2_2
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18353_ rbzero.wall_tracer.trackDistY\[7\] rbzero.wall_tracer.stepDistY\[7\] vssd1
+ vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__or2_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15565_ _08177_ _08178_ vssd1 vssd1 vccd1 vccd1 _08179_ sky130_fd_sc_hd__or2_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12777_ _05459_ _05445_ _05465_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__a21o_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17304_ _09840_ _09842_ vssd1 vssd1 vccd1 vccd1 _09843_ sky130_fd_sc_hd__xor2_1
XFILLER_202_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14516_ _05602_ _07083_ _07140_ _07177_ vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__o2bb2a_2
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18284_ _02046_ _02049_ _02047_ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__o21ai_1
XFILLER_124_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ _04099_ _04409_ _04443_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__nand3b_2
XFILLER_226_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15496_ _08035_ _08109_ vssd1 vssd1 vccd1 vccd1 _08110_ sky130_fd_sc_hd__nand2_1
XFILLER_175_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17235_ _09651_ _09755_ vssd1 vssd1 vccd1 vccd1 _09774_ sky130_fd_sc_hd__nand2_1
XFILLER_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14447_ _05577_ _07124_ _07134_ vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__a21bo_1
XFILLER_70_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11659_ rbzero.tex_g1\[27\] rbzero.tex_g1\[26\] _04374_ vssd1 vssd1 vccd1 vccd1 _04375_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17166_ _08241_ _08917_ vssd1 vssd1 vccd1 vccd1 _09706_ sky130_fd_sc_hd__nor2_1
XFILLER_31_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14378_ _05586_ _07035_ _07066_ vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__o21ai_1
XFILLER_122_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16117_ _08672_ _08674_ _08669_ vssd1 vssd1 vccd1 vccd1 _08729_ sky130_fd_sc_hd__a21bo_1
XFILLER_183_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13329_ _05996_ _06016_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__or2b_1
X_17097_ _09636_ _09637_ vssd1 vssd1 vccd1 vccd1 _09638_ sky130_fd_sc_hd__and2b_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16048_ _08505_ _08522_ _08660_ vssd1 vssd1 vccd1 vccd1 _08661_ sky130_fd_sc_hd__a21bo_1
XFILLER_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19807_ _04111_ _03102_ _03104_ vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__a21oi_1
XFILLER_57_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17999_ _01630_ _01633_ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__nand2_1
XFILLER_111_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19738_ rbzero.pov.ready_buffer\[32\] _03069_ _03070_ rbzero.debug_overlay.facingY\[10\]
+ _03065_ vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__o221a_1
XFILLER_211_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19669_ _07558_ _02836_ _03012_ _03029_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__o211ai_1
XFILLER_225_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20513_ net127 _00529_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20444_ net138 _00475_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20375_ net126 _00406_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10961_ _03708_ vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12700_ _05381_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__inv_2
XFILLER_232_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13680_ _06366_ _06323_ _06364_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__or3_1
XFILLER_243_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10892_ _03672_ vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12631_ _05305_ _05284_ _05316_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__a21o_1
XFILLER_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15350_ _04936_ _07392_ _07393_ _07397_ vssd1 vssd1 vccd1 vccd1 _07964_ sky130_fd_sc_hd__o31a_2
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12562_ rbzero.wall_tracer.rayAddendX\[-2\] _05250_ _05219_ vssd1 vssd1 vccd1 vccd1
+ _05251_ sky130_fd_sc_hd__mux2_2
XFILLER_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14301_ _05531_ vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__buf_2
XFILLER_211_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11513_ _04212_ _04208_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__nor2_1
XFILLER_8_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15281_ _07485_ _07805_ _07802_ _07799_ vssd1 vssd1 vccd1 vccd1 _07895_ sky130_fd_sc_hd__o31a_1
XFILLER_184_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12493_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[10\] vssd1
+ vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__xnor2_2
XFILLER_71_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17020_ _09559_ _09560_ vssd1 vssd1 vccd1 vccd1 _09561_ sky130_fd_sc_hd__nor2_1
XFILLER_172_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14232_ _06735_ _06920_ vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__and2_1
XFILLER_138_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11444_ rbzero.tex_r1\[23\] rbzero.tex_r1\[22\] _04148_ vssd1 vssd1 vccd1 vccd1 _04162_
+ sky130_fd_sc_hd__mux2_1
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14163_ _06829_ _06830_ vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__nor2_1
XFILLER_193_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11375_ _03784_ _04075_ _04072_ _03290_ _04093_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__o221a_1
XFILLER_153_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13114_ _05625_ _05609_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__nor2_1
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10326_ rbzero.tex_r1\[61\] rbzero.tex_r1\[62\] _03366_ vssd1 vssd1 vccd1 vccd1 _03373_
+ sky130_fd_sc_hd__mux2_1
X_14094_ _06707_ _06731_ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__or2_1
XFILLER_193_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18971_ _02645_ vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__clkbuf_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17922_ _01702_ _01704_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__xnor2_1
X_13045_ _05721_ _05733_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__xnor2_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10257_ rbzero.tex_b1\[30\] rbzero.tex_b1\[31\] _03333_ vssd1 vssd1 vccd1 vccd1 _03337_
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17853_ _08240_ _09976_ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__or2_1
XFILLER_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10188_ rbzero.tex_b1\[63\] net50 _03300_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__mux2_1
XFILLER_94_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16804_ _09346_ _09347_ _09348_ vssd1 vssd1 vccd1 vccd1 _09349_ sky130_fd_sc_hd__and3_1
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17784_ _08067_ _08595_ _08645_ _09197_ vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__or4_1
X_14996_ _07606_ _07608_ _07609_ vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__and3_1
XFILLER_82_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19523_ rbzero.pov.spi_buffer\[57\] rbzero.pov.spi_buffer\[58\] _02921_ vssd1 vssd1
+ vccd1 vccd1 _02930_ sky130_fd_sc_hd__mux2_1
XFILLER_75_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13947_ _06579_ _06635_ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__nor2_1
X_16735_ rbzero.wall_tracer.trackDistX\[-11\] rbzero.wall_tracer.stepDistX\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _09288_ sky130_fd_sc_hd__nand2_1
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16666_ rbzero.row_render.size\[3\] _09255_ _07185_ _09259_ vssd1 vssd1 vccd1 vccd1
+ _00501_ sky130_fd_sc_hd__a22o_1
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19454_ rbzero.pov.spi_buffer\[24\] rbzero.pov.spi_buffer\[25\] _02888_ vssd1 vssd1
+ vccd1 vccd1 _02894_ sky130_fd_sc_hd__mux2_1
X_13878_ _06564_ _06566_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__and2_1
XFILLER_34_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15617_ _08228_ _08230_ vssd1 vssd1 vccd1 vccd1 _08231_ sky130_fd_sc_hd__nor2_1
X_18405_ rbzero.debug_overlay.vplaneX\[-9\] _02157_ _02158_ rbzero.wall_tracer.rayAddendX\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a22o_1
XFILLER_201_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12829_ _05497_ _05455_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__nand2_1
X_16597_ _09204_ _09205_ vssd1 vssd1 vccd1 vccd1 _09206_ sky130_fd_sc_hd__nor2_1
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19385_ _02861_ vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__clkinv_2
XFILLER_222_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18336_ _02095_ _02096_ _02097_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__o21a_1
X_15548_ _08150_ _08151_ vssd1 vssd1 vccd1 vccd1 _08162_ sky130_fd_sc_hd__or2b_1
XFILLER_241_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18267_ _01995_ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__clkbuf_4
XFILLER_148_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15479_ _08079_ _08092_ vssd1 vssd1 vccd1 vccd1 _08093_ sky130_fd_sc_hd__xnor2_2
XFILLER_50_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17218_ _09649_ _09650_ _09756_ vssd1 vssd1 vccd1 vccd1 _09758_ sky130_fd_sc_hd__and3_1
XFILLER_200_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18198_ _01894_ _01898_ vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__nand2_1
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17149_ _09687_ _09688_ vssd1 vssd1 vccd1 vccd1 _09689_ sky130_fd_sc_hd__and2b_1
XFILLER_190_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20160_ _03184_ _03185_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__nor2_1
XFILLER_239_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20091_ _03131_ vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__clkinv_2
XFILLER_112_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20993_ net72 _01009_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20427_ net117 _00458_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11160_ _03834_ _03872_ _03878_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__o21ba_2
XFILLER_162_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20358_ gpout3.clk_div\[0\] _03003_ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__nor2_1
XTAP_6202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11091_ _03802_ _03807_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__or2_2
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20289_ _03257_ vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__clkinv_2
XTAP_6246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14850_ _07364_ _07463_ vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__nand2_1
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ _06420_ _06429_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__and2_1
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14781_ rbzero.debug_overlay.playerX\[-5\] _07365_ vssd1 vssd1 vccd1 vccd1 _07395_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_112_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11993_ gpout2.clk_div\[0\] _04664_ net15 vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__and3_1
XFILLER_99_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16520_ _08510_ _08985_ vssd1 vssd1 vccd1 vccd1 _09129_ sky130_fd_sc_hd__nor2_1
XFILLER_21_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13732_ _06166_ _06174_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__nand2_1
X_10944_ _03699_ vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16451_ _08929_ _08930_ vssd1 vssd1 vccd1 vccd1 _09061_ sky130_fd_sc_hd__nand2_1
XFILLER_232_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13663_ _06313_ _06306_ _06309_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__o21a_1
XFILLER_147_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10875_ _03663_ vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15402_ _07973_ _08015_ vssd1 vssd1 vccd1 vccd1 _08016_ sky130_fd_sc_hd__xnor2_2
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ _05220_ _05302_ _05280_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__a21o_1
X_19170_ rbzero.color_sky\[4\] _02752_ _02760_ vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__a21o_1
X_16382_ _08989_ _08990_ vssd1 vssd1 vccd1 vccd1 _08992_ sky130_fd_sc_hd__and2_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13594_ _06280_ _06282_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__xnor2_1
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18121_ _01798_ _01800_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__nor2_1
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15333_ _07933_ _07946_ vssd1 vssd1 vccd1 vccd1 _07947_ sky130_fd_sc_hd__xor2_1
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12545_ _05148_ _05153_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__nor2_1
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18052_ _01832_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__inv_2
X_15264_ _07792_ vssd1 vssd1 vccd1 vccd1 _07878_ sky130_fd_sc_hd__clkbuf_4
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12476_ rbzero.debug_overlay.facingX\[-4\] rbzero.wall_tracer.rayAddendX\[4\] vssd1
+ vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__nor2_1
X_17003_ _09542_ _09543_ vssd1 vssd1 vccd1 vccd1 _09544_ sky130_fd_sc_hd__nor2_1
X_14215_ _06886_ _06902_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__and2_1
X_11427_ _04144_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__buf_2
XANTENNA_5 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ _07807_ _07808_ vssd1 vssd1 vccd1 vccd1 _07809_ sky130_fd_sc_hd__and2b_1
XFILLER_193_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14146_ _06796_ _06797_ _06834_ vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__nand3_1
XFILLER_126_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11358_ _04045_ _04076_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__nand2_1
XFILLER_141_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10309_ rbzero.tex_b1\[5\] rbzero.tex_b1\[6\] _03355_ vssd1 vssd1 vccd1 vccd1 _03364_
+ sky130_fd_sc_hd__mux2_1
XFILLER_193_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14077_ _06470_ _06342_ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__or2_1
X_18954_ _02636_ vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__clkbuf_1
XFILLER_234_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11289_ rbzero.tex_r0\[15\] rbzero.tex_r0\[14\] _03961_ vssd1 vssd1 vccd1 vccd1 _04008_
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17905_ _01685_ _01687_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__nor2_1
X_13028_ _05714_ _05716_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18885_ rbzero.spi_registers.spi_counter\[3\] _02594_ vssd1 vssd1 vccd1 vccd1 _02597_
+ sky130_fd_sc_hd__nand2_1
XTAP_6780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17836_ _10121_ _01589_ _01591_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__a21o_1
XFILLER_227_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17767_ _07618_ _09955_ _10095_ _08732_ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__o22ai_1
XFILLER_130_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14979_ _07592_ vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__buf_2
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19506_ _02865_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__clkbuf_4
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16718_ _04939_ _07254_ rbzero.wall_tracer.state\[1\] vssd1 vssd1 vccd1 vccd1 _09272_
+ sky130_fd_sc_hd__mux2_1
XFILLER_235_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17698_ _01480_ _01481_ _10120_ _10122_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__o211a_1
XFILLER_169_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19437_ rbzero.pov.spi_buffer\[16\] rbzero.pov.spi_buffer\[17\] _02877_ vssd1 vssd1
+ vccd1 vccd1 _02885_ sky130_fd_sc_hd__mux2_1
XFILLER_90_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16649_ _09247_ _03813_ _04228_ vssd1 vssd1 vccd1 vccd1 _09250_ sky130_fd_sc_hd__and3_1
XFILLER_195_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19368_ _02859_ vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__clkinv_2
XFILLER_176_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18319_ _02076_ _02079_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__nand2_1
XFILLER_163_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19299_ _02835_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__buf_2
XFILLER_148_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21330_ _00353_ _01346_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21261_ _00310_ _01277_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20212_ rbzero.traced_texa\[7\] rbzero.texV\[7\] vssd1 vssd1 vccd1 vccd1 _03231_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_117_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21192_ _00241_ _01208_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20143_ _03171_ _03172_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__and2b_1
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20074_ _03130_ vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__clkinv_2
XFILLER_58_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20976_ net63 _00992_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10660_ _03550_ vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10591_ _03514_ vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12330_ _05010_ _04988_ _05017_ _05023_ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__or4_1
XFILLER_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12261_ rbzero.wall_tracer.trackDistX\[-1\] _04953_ rbzero.wall_tracer.trackDistX\[-2\]
+ _04954_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__o22a_1
XFILLER_181_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14000_ _06686_ _06688_ vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__and2b_1
XFILLER_120_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11212_ _03926_ _03927_ _03930_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__mux2_1
X_12192_ _04873_ net35 _04895_ _04897_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__and4_1
XFILLER_122_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11143_ _03846_ _03861_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__or2_1
XTAP_6021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15951_ _07344_ _08564_ vssd1 vssd1 vccd1 vccd1 _08565_ sky130_fd_sc_hd__or2b_1
X_11074_ _03797_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__buf_6
XFILLER_7_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14902_ _04928_ _07515_ vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__nand2_2
XFILLER_231_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15882_ _08493_ _08494_ _08495_ vssd1 vssd1 vccd1 vccd1 _08496_ sky130_fd_sc_hd__nand3_1
XTAP_5364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18670_ _02398_ _02399_ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__or2b_1
XTAP_5375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17621_ _10155_ _10156_ vssd1 vssd1 vccd1 vccd1 _10157_ sky130_fd_sc_hd__nand2_1
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14833_ _07100_ _07204_ _07205_ vssd1 vssd1 vccd1 vccd1 _07447_ sky130_fd_sc_hd__and3_1
XFILLER_40_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ _10087_ _10088_ vssd1 vssd1 vccd1 vccd1 _10089_ sky130_fd_sc_hd__nand2_1
X_14764_ _07377_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__buf_2
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _04665_ _04447_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__nand2_1
XFILLER_229_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16503_ _08982_ _08993_ _09111_ vssd1 vssd1 vccd1 vccd1 _09112_ sky130_fd_sc_hd__a21oi_1
X_13715_ _06398_ _06403_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__or2_1
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17483_ _09757_ _09884_ _09883_ vssd1 vssd1 vccd1 vccd1 _10021_ sky130_fd_sc_hd__a21o_1
XFILLER_32_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10927_ _03690_ vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14695_ rbzero.wall_tracer.stepDistX\[2\] _07208_ _07316_ vssd1 vssd1 vccd1 vccd1
+ _07322_ sky130_fd_sc_hd__mux2_1
XFILLER_60_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19222_ _02792_ vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16434_ _09036_ _09042_ vssd1 vssd1 vccd1 vccd1 _09044_ sky130_fd_sc_hd__or2_1
X_13646_ _06332_ _06334_ _06319_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__a21boi_1
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10858_ _03654_ vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _08862_ _08876_ _08874_ vssd1 vssd1 vccd1 vccd1 _08975_ sky130_fd_sc_hd__a21o_1
XFILLER_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19153_ rbzero.spi_registers.new_leak\[4\] _02745_ vssd1 vssd1 vccd1 vccd1 _02750_
+ sky130_fd_sc_hd__or2_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ _05610_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__clkbuf_4
X_10789_ _03618_ vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__clkbuf_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18104_ _01882_ _01884_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__xor2_1
X_15316_ _07928_ _07929_ vssd1 vssd1 vccd1 vccd1 _07930_ sky130_fd_sc_hd__nand2_1
XFILLER_185_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12528_ rbzero.wall_tracer.visualWallDist\[-1\] _05189_ rbzero.wall_tracer.rcp_sel\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__a21o_1
X_16296_ _08772_ _08905_ _08906_ vssd1 vssd1 vccd1 vccd1 _08907_ sky130_fd_sc_hd__a21oi_1
XFILLER_185_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19084_ _02705_ vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18035_ _01814_ _01816_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__xnor2_1
X_15247_ _07700_ _07860_ _07699_ vssd1 vssd1 vccd1 vccd1 _07861_ sky130_fd_sc_hd__o21ba_1
XFILLER_172_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12459_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__nor2_1
XFILLER_173_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15178_ _07789_ vssd1 vssd1 vccd1 vccd1 _07792_ sky130_fd_sc_hd__buf_2
XFILLER_160_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14129_ _06101_ _06422_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__nor2_1
XFILLER_193_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19986_ _03121_ vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__clkinv_2
XFILLER_154_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18937_ _02627_ vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18868_ rbzero.spi_registers.spi_counter\[1\] _02582_ vssd1 vssd1 vccd1 vccd1 _02583_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_95_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17819_ _01524_ _01602_ vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18799_ _02472_ _04260_ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__or2_1
XFILLER_243_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20830_ _00048_ _00846_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20761_ net107 _00777_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20692_ net70 _00708_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[72\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21313_ net111 _01329_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21244_ _00293_ _01260_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21175_ _00224_ _01191_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20126_ rbzero.traced_texa\[-7\] rbzero.texV\[-7\] vssd1 vssd1 vccd1 vccd1 _03159_
+ sky130_fd_sc_hd__nand2_1
XFILLER_137_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20057_ _03128_ vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__clkinv_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _03902_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__clkbuf_4
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11761_ rbzero.tex_b0\[35\] _04142_ _04144_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__and3_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20959_ net91 _00975_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_202_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13500_ _06187_ _06188_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__nor2_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ rbzero.tex_g1\[8\] rbzero.tex_g1\[9\] _03574_ vssd1 vssd1 vccd1 vccd1 _03578_
+ sky130_fd_sc_hd__mux2_1
X_14480_ _07102_ _07164_ vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__nand2_2
XFILLER_42_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _03900_ _04395_ _04399_ _03985_ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__o311a_1
XFILLER_241_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _06114_ _06118_ _06119_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__nor3_1
XFILLER_186_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10643_ rbzero.tex_g1\[41\] rbzero.tex_g1\[42\] _03541_ vssd1 vssd1 vccd1 vccd1 _03542_
+ sky130_fd_sc_hd__mux2_1
XFILLER_224_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16150_ _08759_ _08761_ vssd1 vssd1 vccd1 vccd1 _08762_ sky130_fd_sc_hd__xor2_1
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13362_ _05607_ _06050_ _06008_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__mux2_1
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10574_ _03505_ vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__clkbuf_1
X_15101_ _07683_ _07714_ vssd1 vssd1 vccd1 vccd1 _07715_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12313_ rbzero.wall_tracer.trackDistX\[6\] _05004_ rbzero.wall_tracer.trackDistX\[5\]
+ _05002_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__a22o_1
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16081_ _08553_ _08554_ vssd1 vssd1 vccd1 vccd1 _08694_ sky130_fd_sc_hd__or2_1
XFILLER_154_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13293_ _05942_ _05944_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15032_ _07645_ vssd1 vssd1 vccd1 vccd1 _07646_ sky130_fd_sc_hd__clkbuf_4
XFILLER_170_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12244_ _04937_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__buf_4
XFILLER_108_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19840_ _03107_ vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__clkinv_2
XFILLER_155_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12175_ _04871_ _04880_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__or2_1
XFILLER_68_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11126_ rbzero.texV\[4\] _03843_ _03844_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__a21boi_1
X_19771_ _03289_ _03443_ _03803_ _03078_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__or4_1
X_16983_ _09420_ _09517_ _09522_ vssd1 vssd1 vccd1 vccd1 _09524_ sky130_fd_sc_hd__and3_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18722_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.debug_overlay.vplaneY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__or2_1
X_15934_ _07900_ _08530_ _08547_ vssd1 vssd1 vccd1 vccd1 _08548_ sky130_fd_sc_hd__a21o_1
XTAP_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11057_ _03783_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__clkbuf_4
XFILLER_237_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18653_ rbzero.debug_overlay.vplaneY\[-9\] _02166_ _02158_ rbzero.wall_tracer.rayAddendY\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__a22o_1
X_15865_ _07470_ _07471_ _07834_ _08478_ vssd1 vssd1 vccd1 vccd1 _08479_ sky130_fd_sc_hd__or4_1
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17604_ _10139_ _10140_ vssd1 vssd1 vccd1 vccd1 _10141_ sky130_fd_sc_hd__xnor2_1
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14816_ rbzero.wall_tracer.visualWallDist\[-8\] _03793_ rbzero.wall_tracer.state\[6\]
+ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__a21oi_1
X_18584_ _02324_ vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__clkbuf_1
X_15796_ _08404_ _08406_ _08409_ vssd1 vssd1 vccd1 vccd1 _08410_ sky130_fd_sc_hd__o21ai_1
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17535_ _09957_ _09959_ _09956_ vssd1 vssd1 vccd1 vccd1 _10072_ sky130_fd_sc_hd__a21bo_1
XFILLER_166_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_143 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_143/HI o_rgb[1] sky130_fd_sc_hd__conb_1
XFILLER_79_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14747_ _07339_ _05113_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__nand2_1
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11959_ _04664_ _04665_ _04668_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__or3_1
Xtop_ew_algofoogle_154 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_154/HI o_rgb[16]
+ sky130_fd_sc_hd__conb_1
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17466_ _10001_ _10003_ vssd1 vssd1 vccd1 vccd1 _10004_ sky130_fd_sc_hd__xor2_1
X_14678_ rbzero.wall_tracer.stepDistX\[-6\] _07180_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _07313_ sky130_fd_sc_hd__mux2_1
XFILLER_220_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19205_ rbzero.spi_registers.vshift\[5\] _02774_ _02782_ _02780_ vssd1 vssd1 vccd1
+ vccd1 _00766_ sky130_fd_sc_hd__o211a_1
X_16417_ _09025_ _09026_ vssd1 vssd1 vccd1 vccd1 _09027_ sky130_fd_sc_hd__nand2_1
X_13629_ _05818_ _06306_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__nand2_1
XFILLER_203_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17397_ _09833_ _07619_ _09571_ _08671_ vssd1 vssd1 vccd1 vccd1 _09935_ sky130_fd_sc_hd__o22ai_1
XFILLER_34_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19136_ rbzero.othery\[4\] _02723_ _02737_ _02738_ vssd1 vssd1 vccd1 vccd1 _00741_
+ sky130_fd_sc_hd__o211a_1
XFILLER_203_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16348_ _08839_ _08958_ vssd1 vssd1 vccd1 vccd1 _08959_ sky130_fd_sc_hd__xor2_4
XFILLER_158_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16279_ _08274_ vssd1 vssd1 vccd1 vccd1 _08890_ sky130_fd_sc_hd__buf_2
XFILLER_12_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19067_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.spi_buffer\[4\]
+ _02690_ vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__mux2_1
XFILLER_195_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18018_ _01648_ _01684_ _01799_ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__a21oi_1
XFILLER_195_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout106 net108 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_2
Xfanout117 net122 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout128 net129 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_2
XFILLER_134_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout139 net140 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_4
XFILLER_141_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19969_ _03119_ vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__clkinv_2
XFILLER_234_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20813_ _00031_ _00829_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20744_ net105 _00760_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20675_ net68 _00691_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10290_ rbzero.tex_b1\[14\] rbzero.tex_b1\[15\] _03344_ vssd1 vssd1 vccd1 vccd1 _03354_
+ sky130_fd_sc_hd__mux2_1
XFILLER_191_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21227_ _00276_ _01243_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21158_ _00207_ _01174_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20109_ rbzero.traced_texa\[-10\] rbzero.texV\[-10\] vssd1 vssd1 vccd1 vccd1 _03145_
+ sky130_fd_sc_hd__nand2_1
XFILLER_8_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13980_ _06470_ _06330_ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__nor2_1
X_21089_ _00138_ _01105_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12931_ _05607_ _05610_ _05619_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__or3_1
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12862_ _05481_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__or2_1
X_15650_ _08196_ _08206_ vssd1 vssd1 vccd1 vccd1 _08264_ sky130_fd_sc_hd__xnor2_1
XFILLER_160_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _04965_ _07246_ _07249_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__o21ai_1
X_11813_ rbzero.tex_b1\[63\] rbzero.tex_b1\[62\] _04032_ vssd1 vssd1 vccd1 vccd1 _04527_
+ sky130_fd_sc_hd__mux2_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _08176_ _08175_ vssd1 vssd1 vccd1 vccd1 _08195_ sky130_fd_sc_hd__and2_1
XFILLER_160_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12793_ _05480_ _05481_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__nor2_1
XFILLER_15_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _09733_ _09735_ _09858_ vssd1 vssd1 vccd1 vccd1 _09859_ sky130_fd_sc_hd__nand3_1
XFILLER_242_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14532_ _07207_ vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11744_ rbzero.tex_b0\[54\] _03959_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__and2_1
XFILLER_202_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17251_ _09699_ _09715_ vssd1 vssd1 vccd1 vccd1 _09790_ sky130_fd_sc_hd__or2b_1
X_14463_ _06987_ _07030_ _07121_ _05517_ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__a22oi_1
XFILLER_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11675_ _03994_ _04386_ _04390_ _03900_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__a211o_1
XFILLER_174_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16202_ _08746_ _08813_ vssd1 vssd1 vccd1 vccd1 _08814_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13414_ _05699_ _05641_ _05651_ _05612_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__a22o_1
XFILLER_146_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17182_ _08787_ _09207_ _09449_ vssd1 vssd1 vccd1 vccd1 _09722_ sky130_fd_sc_hd__a21o_1
XFILLER_179_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10626_ rbzero.tex_g1\[49\] rbzero.tex_g1\[50\] _03530_ vssd1 vssd1 vccd1 vccd1 _03533_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14394_ _07007_ _07082_ _07079_ _07025_ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16133_ _08715_ _08744_ vssd1 vssd1 vccd1 vccd1 _08745_ sky130_fd_sc_hd__xnor2_1
X_13345_ _05793_ _05749_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__nor2_1
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10557_ _03496_ vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16064_ _08675_ _08676_ vssd1 vssd1 vccd1 vccd1 _08677_ sky130_fd_sc_hd__and2b_1
XFILLER_182_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13276_ _05963_ _05964_ _05635_ _05638_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__a211o_1
XFILLER_127_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10488_ _03460_ vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15015_ _07518_ _07530_ _07627_ vssd1 vssd1 vccd1 vccd1 _07629_ sky130_fd_sc_hd__nand3_1
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12227_ _03817_ _03730_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__nor2_1
XFILLER_194_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19823_ _03105_ vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__clkinv_2
XFILLER_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12158_ _04825_ net27 gpout4.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__and3_1
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11109_ rbzero.traced_texVinit\[6\] rbzero.spi_registers.vshift\[3\] vssd1 vssd1
+ vccd1 vccd1 _03828_ sky130_fd_sc_hd__or2_1
XFILLER_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19754_ rbzero.pov.ready_buffer\[4\] _03055_ _03058_ rbzero.debug_overlay.vplaneY\[-5\]
+ _02832_ vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__o221a_1
X_16966_ _09351_ _09507_ vssd1 vssd1 vccd1 vccd1 _09508_ sky130_fd_sc_hd__nand2_1
X_12089_ net25 net26 vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__and2b_1
XFILLER_231_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18705_ _02427_ _02431_ _03818_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__o21ai_1
X_15917_ rbzero.wall_tracer.visualWallDist\[6\] _03796_ vssd1 vssd1 vccd1 vccd1 _08531_
+ sky130_fd_sc_hd__nand2_4
XFILLER_110_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19685_ rbzero.debug_overlay.playerY\[2\] _03016_ _03042_ _03031_ vssd1 vssd1 vccd1
+ vccd1 _00986_ sky130_fd_sc_hd__o211a_1
X_16897_ _07751_ _07834_ _09170_ vssd1 vssd1 vccd1 vccd1 _09439_ sky130_fd_sc_hd__or3_1
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18636_ rbzero.debug_overlay.playerX\[4\] _02368_ _03797_ vssd1 vssd1 vccd1 vccd1
+ _02369_ sky130_fd_sc_hd__mux2_1
X_15848_ _07815_ _07828_ _07825_ vssd1 vssd1 vccd1 vccd1 _08462_ sky130_fd_sc_hd__a21boi_1
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18567_ _02307_ _02308_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__nand2_1
XFILLER_240_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15779_ _07616_ _07675_ vssd1 vssd1 vccd1 vccd1 _08393_ sky130_fd_sc_hd__nor2_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17518_ _10053_ _10054_ vssd1 vssd1 vccd1 vccd1 _10055_ sky130_fd_sc_hd__xnor2_1
XFILLER_233_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18498_ rbzero.wall_tracer.rayAddendX\[2\] _00013_ _02244_ vssd1 vssd1 vccd1 vccd1
+ _00597_ sky130_fd_sc_hd__o21a_1
XFILLER_221_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17449_ _07814_ _09976_ vssd1 vssd1 vccd1 vccd1 _09987_ sky130_fd_sc_hd__nor2_1
XFILLER_178_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20460_ net126 _00010_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[13\] sky130_fd_sc_hd__dfxtp_2
XFILLER_158_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19119_ rbzero.otherx\[1\] _02723_ _02729_ _02728_ vssd1 vssd1 vccd1 vccd1 _00733_
+ sky130_fd_sc_hd__o211a_1
XFILLER_203_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20391_ net135 _00422_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21012_ net80 _01028_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_102_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20727_ net100 _00743_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11460_ rbzero.tex_r1\[9\] rbzero.tex_r1\[8\] _04168_ vssd1 vssd1 vccd1 vccd1 _04178_
+ sky130_fd_sc_hd__mux2_1
X_20658_ net63 _00674_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10411_ rbzero.tex_r1\[21\] rbzero.tex_r1\[22\] _03411_ vssd1 vssd1 vccd1 vccd1 _03418_
+ sky130_fd_sc_hd__mux2_1
XFILLER_178_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11391_ gpout0.vpos\[9\] vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__buf_2
X_20589_ net95 _00605_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13130_ _05699_ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__nand2_1
XFILLER_125_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10342_ _03381_ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13061_ _05608_ _05749_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__nor2_1
XFILLER_69_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10273_ _03345_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12012_ _04719_ _04720_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__nand2_1
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16820_ rbzero.wall_tracer.trackDistX\[-1\] rbzero.wall_tracer.stepDistX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _09363_ sky130_fd_sc_hd__and2_1
XFILLER_120_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16751_ _07332_ _08576_ vssd1 vssd1 vccd1 vccd1 _09302_ sky130_fd_sc_hd__and2_1
X_13963_ _06594_ _06651_ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__nor2_1
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15702_ _08245_ _08269_ vssd1 vssd1 vccd1 vccd1 _08316_ sky130_fd_sc_hd__nor2_1
XFILLER_235_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12914_ _05568_ _05598_ _05601_ _05602_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__o31a_1
X_19470_ _02902_ vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__clkbuf_1
XFILLER_234_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13894_ _06577_ _06582_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__or2_1
X_16682_ _09254_ vssd1 vssd1 vccd1 vccd1 _09262_ sky130_fd_sc_hd__clkbuf_4
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18421_ rbzero.debug_overlay.vplaneX\[-3\] rbzero.wall_tracer.rayAddendX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__nand2_1
X_15633_ _08244_ _08246_ vssd1 vssd1 vccd1 vccd1 _08247_ sky130_fd_sc_hd__and2b_1
X_12845_ _05478_ _05454_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__or2_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ rbzero.wall_tracer.trackDistY\[6\] _02039_ _02112_ _01506_ vssd1 vssd1 vccd1
+ vccd1 _00583_ sky130_fd_sc_hd__o22a_1
XFILLER_37_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _08117_ _08120_ vssd1 vssd1 vccd1 vccd1 _08178_ sky130_fd_sc_hd__xnor2_1
X_12776_ _05417_ _05438_ _05350_ _05372_ _05448_ _05444_ vssd1 vssd1 vccd1 vccd1 _05465_
+ sky130_fd_sc_hd__mux4_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _08760_ _08628_ _09708_ _09841_ vssd1 vssd1 vccd1 vccd1 _09842_ sky130_fd_sc_hd__o31a_1
XFILLER_163_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ _07194_ vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11727_ _03954_ _04417_ _04425_ _04442_ _03896_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__a311o_1
X_18283_ rbzero.wall_tracer.trackDistY\[-3\] rbzero.wall_tracer.stepDistY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__nand2_1
X_15495_ _08036_ _08108_ vssd1 vssd1 vccd1 vccd1 _08109_ sky130_fd_sc_hd__or2_1
XFILLER_148_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17234_ _09752_ _09754_ vssd1 vssd1 vccd1 vccd1 _09773_ sky130_fd_sc_hd__or2_1
XFILLER_204_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14446_ _05577_ _07129_ _07132_ _07133_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__o31a_1
XFILLER_128_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11658_ _03974_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__clkbuf_4
XFILLER_122_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10609_ rbzero.tex_g1\[57\] rbzero.tex_g1\[58\] _03519_ vssd1 vssd1 vccd1 vccd1 _03524_
+ sky130_fd_sc_hd__mux2_1
X_17165_ _09703_ _09704_ vssd1 vssd1 vccd1 vccd1 _09705_ sky130_fd_sc_hd__xor2_1
X_14377_ _05501_ _07042_ _07043_ vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__or3_1
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11589_ rbzero.tex_g0\[21\] rbzero.tex_g0\[20\] _04119_ vssd1 vssd1 vccd1 vccd1 _04306_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16116_ _08664_ _08727_ vssd1 vssd1 vccd1 vccd1 _08728_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13328_ _05996_ _06016_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17096_ _09514_ _09515_ _09635_ vssd1 vssd1 vccd1 vccd1 _09637_ sky130_fd_sc_hd__a21o_1
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16047_ _08523_ _08503_ vssd1 vssd1 vccd1 vccd1 _08660_ sky130_fd_sc_hd__or2b_1
XFILLER_170_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13259_ _05938_ _05947_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__and2b_1
XFILLER_171_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19806_ _04110_ _03808_ _03103_ _02708_ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__a31o_1
XFILLER_233_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17998_ _01671_ _01672_ _01674_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__a21bo_1
XFILLER_96_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19737_ _03058_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__clkbuf_4
X_16949_ _09181_ _09219_ _09490_ vssd1 vssd1 vccd1 vccd1 _09491_ sky130_fd_sc_hd__a21o_1
XFILLER_226_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19668_ rbzero.pov.ready_buffer\[52\] _02836_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__nand2_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18619_ _03735_ _07491_ _02349_ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__o21ai_1
XFILLER_213_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19599_ rbzero.pov.ready_buffer\[66\] _07546_ _02962_ vssd1 vssd1 vccd1 vccd1 _02976_
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20512_ net127 _00528_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20443_ net137 _00474_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20374_ net118 _00012_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rcp_sel\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10960_ rbzero.tex_b0\[19\] rbzero.tex_b0\[18\] _03704_ vssd1 vssd1 vccd1 vccd1 _03708_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10891_ rbzero.tex_b0\[52\] rbzero.tex_b0\[51\] _03671_ vssd1 vssd1 vccd1 vccd1 _03672_
+ sky130_fd_sc_hd__mux2_1
XFILLER_232_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12630_ _05187_ _05288_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__nand2_1
XFILLER_245_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12561_ rbzero.wall_tracer.visualWallDist\[-10\] rbzero.wall_tracer.rayAddendY\[-2\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__mux2_1
XFILLER_93_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14300_ _05434_ _06987_ _06988_ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__or3b_1
XFILLER_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ _04222_ _04227_ _04229_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__o21ba_1
XFILLER_200_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15280_ _07892_ _07893_ vssd1 vssd1 vccd1 vccd1 _07894_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12492_ _05146_ _05177_ _05180_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__o21bai_1
XFILLER_141_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14231_ _06137_ _06172_ vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__nor2_1
XFILLER_71_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11443_ rbzero.tex_r1\[21\] rbzero.tex_r1\[20\] _04000_ vssd1 vssd1 vccd1 vccd1 _04161_
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14162_ _06845_ _06848_ _06850_ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__a21o_1
XFILLER_125_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11374_ _03781_ _04077_ _04075_ _03783_ _04092_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__a221o_1
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13113_ _05786_ _05801_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__xnor2_1
X_10325_ _03372_ vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__clkbuf_1
X_14093_ _06733_ _06781_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__nor2_1
XFILLER_125_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18970_ rbzero.pov.spi_buffer\[33\] rbzero.pov.ready_buffer\[33\] _02640_ vssd1 vssd1
+ vccd1 vccd1 _02645_ sky130_fd_sc_hd__mux2_1
XFILLER_180_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ _01524_ _01602_ _01703_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__a21oi_2
X_13044_ _05724_ _05732_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__xor2_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10256_ _03336_ vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17852_ _01633_ _01634_ vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__and2_1
XFILLER_121_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10187_ _03299_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__clkbuf_4
XTAP_6984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16803_ _09339_ _09342_ _09340_ vssd1 vssd1 vccd1 vccd1 _09348_ sky130_fd_sc_hd__o21ai_1
X_17783_ _01476_ _01478_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__nand2_1
XFILLER_130_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14995_ _07566_ _07593_ vssd1 vssd1 vccd1 vccd1 _07609_ sky130_fd_sc_hd__nor2_1
XFILLER_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19522_ _02929_ vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__clkbuf_1
X_16734_ rbzero.wall_tracer.trackDistX\[-11\] rbzero.wall_tracer.stepDistX\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _09287_ sky130_fd_sc_hd__or2_1
X_13946_ _05767_ _06634_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__or2_1
XFILLER_130_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19453_ _02893_ vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__clkbuf_1
X_16665_ rbzero.row_render.size\[2\] _09255_ _07180_ _09259_ vssd1 vssd1 vccd1 vccd1
+ _00500_ sky130_fd_sc_hd__a22o_1
XFILLER_235_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13877_ _06450_ _06565_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__nor2_1
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18404_ _03810_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__buf_4
XFILLER_179_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15616_ _08180_ _08229_ vssd1 vssd1 vccd1 vccd1 _08230_ sky130_fd_sc_hd__xnor2_1
X_12828_ _05515_ _05516_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__nand2_2
X_19384_ _02861_ vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__clkinv_2
X_16596_ _07826_ _09197_ _09202_ _09203_ vssd1 vssd1 vccd1 vccd1 _09205_ sky130_fd_sc_hd__o22a_1
XFILLER_201_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18335_ _02095_ _02096_ _02097_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__nor3_1
X_15547_ _08115_ _08160_ vssd1 vssd1 vccd1 vccd1 _08161_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12759_ _05428_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__clkbuf_4
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18266_ rbzero.wall_tracer.trackDistY\[-6\] _01996_ _02038_ _09324_ vssd1 vssd1 vccd1
+ vccd1 _00571_ sky130_fd_sc_hd__o22a_1
X_15478_ _08080_ _08090_ _08091_ vssd1 vssd1 vccd1 vccd1 _08092_ sky130_fd_sc_hd__a21o_1
XFILLER_147_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17217_ _09649_ _09650_ _09756_ vssd1 vssd1 vccd1 vccd1 _09757_ sky130_fd_sc_hd__a21o_1
XFILLER_175_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14429_ _07102_ _07117_ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__nand2_1
X_18197_ _01894_ _01898_ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__nor2_1
XFILLER_129_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17148_ _09679_ _09686_ vssd1 vssd1 vccd1 vccd1 _09688_ sky130_fd_sc_hd__or2_1
XFILLER_143_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17079_ _09481_ _09483_ vssd1 vssd1 vccd1 vccd1 _09620_ sky130_fd_sc_hd__or2b_1
XFILLER_89_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20090_ _03131_ vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__clkinv_2
XFILLER_135_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20992_ net65 _01008_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20426_ net117 _00457_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20357_ _03281_ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11090_ _03812_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__buf_4
XTAP_6236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20288_ _03257_ vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__clkinv_2
XTAP_5502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13800_ _06478_ _06488_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__or2_1
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14780_ rbzero.debug_overlay.playerX\[-5\] vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__inv_2
XFILLER_21_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11992_ net107 vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__buf_4
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13731_ _06392_ _06419_ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__nand2_1
X_10943_ rbzero.tex_b0\[27\] rbzero.tex_b0\[26\] _03693_ vssd1 vssd1 vccd1 vccd1 _03699_
+ sky130_fd_sc_hd__mux2_1
XFILLER_244_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16450_ _09056_ _09057_ _09058_ vssd1 vssd1 vccd1 vccd1 _09060_ sky130_fd_sc_hd__a21o_1
X_13662_ _06329_ _06338_ _06350_ vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__o21ai_1
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10874_ rbzero.tex_b0\[60\] rbzero.tex_b0\[59\] _03660_ vssd1 vssd1 vccd1 vccd1 _03663_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15401_ _07468_ _07388_ vssd1 vssd1 vccd1 vccd1 _08015_ sky130_fd_sc_hd__nor2_1
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12613_ _05301_ _03816_ _05188_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__o21ai_1
XFILLER_223_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16381_ _08989_ _08990_ vssd1 vssd1 vccd1 vccd1 _08991_ sky130_fd_sc_hd__nor2_1
X_13593_ _06204_ _06245_ _06281_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__o21bai_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18120_ _01892_ _01900_ vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__xnor2_1
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15332_ _07942_ _07945_ vssd1 vssd1 vccd1 vccd1 _07946_ sky130_fd_sc_hd__and2_1
X_12544_ rbzero.wall_tracer.rcp_sel\[0\] _05230_ _05231_ _05232_ vssd1 vssd1 vccd1
+ vccd1 _05233_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_223_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18051_ _01711_ _01819_ _01831_ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__o21a_1
X_15263_ _07746_ _07754_ vssd1 vssd1 vccd1 vccd1 _07877_ sky130_fd_sc_hd__or2b_1
XFILLER_185_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12475_ _05159_ _05160_ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__and3_1
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17002_ _09540_ _09541_ vssd1 vssd1 vccd1 vccd1 _09543_ sky130_fd_sc_hd__and2_1
XFILLER_201_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14214_ _06886_ _06902_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__nor2_1
X_11426_ _03940_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__clkbuf_4
X_15194_ _07804_ _07806_ vssd1 vssd1 vccd1 vccd1 _07808_ sky130_fd_sc_hd__nand2_1
XFILLER_32_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_6 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14145_ _06811_ _06832_ _06833_ vssd1 vssd1 vccd1 vccd1 _06834_ sky130_fd_sc_hd__a21o_1
X_11357_ rbzero.row_render.size\[4\] _04044_ rbzero.row_render.size\[5\] vssd1 vssd1
+ vccd1 vccd1 _04076_ sky130_fd_sc_hd__o21ai_1
XFILLER_158_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10308_ _03363_ vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__clkbuf_1
X_14076_ _05959_ _06331_ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__nor2_1
X_18953_ rbzero.pov.spi_buffer\[25\] rbzero.pov.ready_buffer\[25\] _02629_ vssd1 vssd1
+ vccd1 vccd1 _02636_ sky130_fd_sc_hd__mux2_1
XFILLER_193_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11288_ _03923_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__buf_4
XFILLER_239_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17904_ _01564_ _01598_ _01686_ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__a21boi_2
X_13027_ _05706_ _05707_ _05715_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__a21oi_1
X_10239_ _03327_ vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18884_ _02596_ vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__clkbuf_1
XTAP_6770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17835_ _01612_ _01618_ rbzero.wall_tracer.trackDistX\[7\] _09276_ vssd1 vssd1 vccd1
+ vccd1 _00560_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_67_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17766_ _07618_ _08732_ _09955_ _10095_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__or4_1
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14978_ _04928_ rbzero.wall_tracer.stepDistX\[-10\] _07521_ vssd1 vssd1 vccd1 vccd1
+ _07592_ sky130_fd_sc_hd__o21ai_4
XFILLER_81_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19505_ _02920_ vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__clkbuf_1
XFILLER_130_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16717_ _09271_ vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13929_ _06607_ _06616_ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__nor2_1
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17697_ _10120_ _10122_ _01480_ _01481_ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__a211oi_1
XFILLER_223_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19436_ _02884_ vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__clkbuf_1
XFILLER_222_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16648_ _04203_ _09244_ vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__nor2_1
XFILLER_126_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19367_ _02859_ vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__clkinv_2
XFILLER_76_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16579_ _08478_ _08928_ _08272_ vssd1 vssd1 vccd1 vccd1 _09188_ sky130_fd_sc_hd__a21o_1
XFILLER_124_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18318_ rbzero.wall_tracer.trackDistY\[2\] rbzero.wall_tracer.stepDistY\[2\] vssd1
+ vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__or2_1
XFILLER_163_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19298_ _02834_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__buf_2
XFILLER_198_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18249_ _02021_ _02022_ _02023_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__or3_1
XFILLER_136_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21260_ _00309_ _01276_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20211_ rbzero.texV\[6\] _03137_ _03142_ _03230_ vssd1 vssd1 vccd1 vccd1 _01324_
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21191_ _00240_ _01207_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20142_ rbzero.traced_texa\[-4\] rbzero.texV\[-4\] vssd1 vssd1 vccd1 vccd1 _03172_
+ sky130_fd_sc_hd__nand2_1
XFILLER_137_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20073_ _03130_ vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__clkinv_2
XFILLER_100_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20975_ net90 _00991_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10590_ rbzero.tex_r0\[3\] rbzero.tex_r0\[2\] _03512_ vssd1 vssd1 vccd1 vccd1 _03514_
+ sky130_fd_sc_hd__mux2_1
XFILLER_224_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12260_ rbzero.wall_tracer.trackDistY\[-2\] vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__inv_2
XFILLER_177_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11211_ _03929_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__buf_4
X_20409_ net130 _00440_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_181_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12191_ _04883_ o_rgb[23] _04896_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__a21bo_1
XFILLER_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21389_ net109 _01405_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11142_ _03842_ _03845_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__and2_1
XFILLER_218_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15950_ _08459_ _08563_ vssd1 vssd1 vccd1 vccd1 _08564_ sky130_fd_sc_hd__xor2_2
X_11073_ rbzero.wall_tracer.state\[1\] vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__buf_6
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14901_ _04932_ _07100_ _07146_ _07514_ vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__a31o_2
XFILLER_76_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15881_ _07830_ _07851_ _07850_ vssd1 vssd1 vccd1 vccd1 _08495_ sky130_fd_sc_hd__a21bo_1
XTAP_5365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17620_ _10065_ _10068_ _10154_ vssd1 vssd1 vccd1 vccd1 _10156_ sky130_fd_sc_hd__nand3_1
XTAP_5387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14832_ _07177_ _07162_ _07201_ _07100_ vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__o211a_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17551_ _10049_ _10050_ _10086_ vssd1 vssd1 vccd1 vccd1 _10088_ sky130_fd_sc_hd__nand3_1
XFILLER_217_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14763_ _07356_ _07362_ _07363_ _07376_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__o31ai_4
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11975_ _04681_ _04683_ _04684_ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__and3_1
XFILLER_189_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16502_ _09110_ _08991_ vssd1 vssd1 vccd1 vccd1 _09111_ sky130_fd_sc_hd__xnor2_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13714_ _06383_ _06397_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__nor2_1
X_17482_ _10018_ _10019_ vssd1 vssd1 vccd1 vccd1 _10020_ sky130_fd_sc_hd__or2_1
XFILLER_204_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10926_ rbzero.tex_b0\[35\] rbzero.tex_b0\[34\] _03682_ vssd1 vssd1 vccd1 vccd1 _03690_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14694_ _07321_ vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19221_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.new_sky\[5\] _02786_
+ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__mux2_1
X_16433_ _09036_ _09042_ vssd1 vssd1 vccd1 vccd1 _09043_ sky130_fd_sc_hd__nand2_1
XFILLER_232_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13645_ _06317_ _06333_ _06318_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__mux2_1
X_10857_ rbzero.tex_g0\[4\] rbzero.tex_g0\[3\] _03649_ vssd1 vssd1 vccd1 vccd1 _03654_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19152_ rbzero.floor_leak\[3\] _02744_ _02749_ _02738_ vssd1 vssd1 vccd1 vccd1 _00746_
+ sky130_fd_sc_hd__o211a_1
X_16364_ _08972_ _08973_ vssd1 vssd1 vccd1 vccd1 _08974_ sky130_fd_sc_hd__nor2_1
XFILLER_201_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13576_ _06229_ _06247_ _06248_ _06264_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__a31o_1
XFILLER_169_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10788_ rbzero.tex_g0\[37\] rbzero.tex_g0\[36\] _03616_ vssd1 vssd1 vccd1 vccd1 _03618_
+ sky130_fd_sc_hd__mux2_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _01780_ _01788_ _01883_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__a21oi_1
XFILLER_201_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15315_ _07906_ _07907_ _07927_ vssd1 vssd1 vccd1 vccd1 _07929_ sky130_fd_sc_hd__a21o_1
XFILLER_173_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12527_ _03815_ _05056_ _05099_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__and3_1
X_19083_ rbzero.spi_registers.spi_cmd\[0\] rbzero.spi_registers.spi_cmd\[1\] _02703_
+ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__mux2_1
X_16295_ _08046_ _08771_ _07837_ _08636_ vssd1 vssd1 vccd1 vccd1 _08906_ sky130_fd_sc_hd__and4_1
XFILLER_200_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18034_ _01518_ _01815_ _01698_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__o21a_1
XFILLER_173_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15246_ _07713_ vssd1 vssd1 vccd1 vccd1 _07860_ sky130_fd_sc_hd__inv_2
XFILLER_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12458_ rbzero.debug_overlay.facingX\[-6\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__nor2_1
XFILLER_160_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11409_ rbzero.tex_r1\[63\] rbzero.tex_r1\[62\] _03935_ vssd1 vssd1 vccd1 vccd1 _04127_
+ sky130_fd_sc_hd__mux2_1
XFILLER_236_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15177_ _07501_ _07789_ _07790_ _07575_ vssd1 vssd1 vccd1 vccd1 _07791_ sky130_fd_sc_hd__or4_1
X_12389_ _05044_ _05043_ _05047_ rbzero.wall_tracer.rayAddendY\[3\] rbzero.debug_overlay.facingY\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__a32o_1
XFILLER_193_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14128_ _06765_ _06768_ vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19985_ _03121_ vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__clkinv_2
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14059_ _06741_ _06747_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__or2_1
XFILLER_140_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18936_ rbzero.pov.spi_buffer\[17\] rbzero.pov.ready_buffer\[17\] _02618_ vssd1 vssd1
+ vccd1 vccd1 _02627_ sky130_fd_sc_hd__mux2_1
XFILLER_234_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18867_ rbzero.spi_registers.spi_cmd\[3\] _02581_ rbzero.spi_registers.spi_cmd\[1\]
+ rbzero.spi_registers.spi_cmd\[0\] vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__and4b_1
XFILLER_228_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17818_ _01599_ _01601_ vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__xor2_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18798_ _02505_ _02513_ _02517_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__a21o_1
XFILLER_236_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17749_ _01531_ _01532_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20760_ net105 _00776_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19419_ _02875_ vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__clkbuf_1
XFILLER_223_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20691_ net70 _00707_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[71\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21312_ net111 _01328_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21243_ _00292_ _01259_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21174_ _00223_ _01190_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20125_ rbzero.traced_texa\[-7\] rbzero.texV\[-7\] vssd1 vssd1 vccd1 vccd1 _03158_
+ sky130_fd_sc_hd__or2_1
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20056_ _03128_ vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__clkinv_2
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11760_ rbzero.tex_b0\[33\] rbzero.tex_b0\[32\] _03904_ vssd1 vssd1 vccd1 vccd1 _04475_
+ sky130_fd_sc_hd__mux2_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20958_ net70 _00974_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _03577_ vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_241_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _04007_ _04402_ _04406_ _03956_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__a211o_1
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20889_ net64 _00905_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_201_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13430_ _06099_ _06100_ _06113_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__a21oi_1
X_10642_ _03388_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__clkbuf_4
XFILLER_220_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13361_ _05634_ _05636_ _05629_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10573_ rbzero.tex_r0\[11\] rbzero.tex_r0\[10\] _03501_ vssd1 vssd1 vccd1 vccd1 _03505_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15100_ _07701_ _07713_ vssd1 vssd1 vccd1 vccd1 _07714_ sky130_fd_sc_hd__xnor2_1
XFILLER_167_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12312_ _05003_ _05005_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__nand2_1
XFILLER_33_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16080_ _08691_ _08692_ vssd1 vssd1 vccd1 vccd1 _08693_ sky130_fd_sc_hd__xnor2_1
X_13292_ _05948_ _05975_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__xnor2_2
XFILLER_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15031_ _07644_ vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__clkbuf_4
X_12243_ _04936_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__buf_4
XFILLER_177_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12174_ _03288_ _04592_ _04631_ _04632_ _04874_ _04876_ vssd1 vssd1 vccd1 vccd1 _04880_
+ sky130_fd_sc_hd__mux4_1
XFILLER_122_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11125_ rbzero.traced_texVinit\[4\] rbzero.spi_registers.vshift\[1\] vssd1 vssd1
+ vccd1 vccd1 _03844_ sky130_fd_sc_hd__nand2_1
X_19770_ _04080_ _04591_ _04592_ _04078_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__or4b_1
XFILLER_110_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16982_ _09420_ _09517_ _09522_ vssd1 vssd1 vccd1 vccd1 _09523_ sky130_fd_sc_hd__a21oi_1
XFILLER_231_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18721_ _02443_ _02444_ _02445_ _02442_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__a22o_1
X_15933_ _08532_ _08546_ vssd1 vssd1 vccd1 vccd1 _08547_ sky130_fd_sc_hd__xnor2_1
XTAP_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11056_ gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__clkbuf_4
XFILLER_114_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18652_ _02371_ _02372_ _02382_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__o21ai_1
XFILLER_97_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15864_ _08473_ _08477_ _04937_ vssd1 vssd1 vccd1 vccd1 _08478_ sky130_fd_sc_hd__a21o_2
XTAP_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17603_ _09912_ _10010_ _10008_ vssd1 vssd1 vccd1 vccd1 _10140_ sky130_fd_sc_hd__a21oi_1
XFILLER_224_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14815_ _07349_ _07428_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__nand2_1
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18583_ rbzero.wall_tracer.rayAddendX\[8\] _02323_ _03812_ vssd1 vssd1 vccd1 vccd1
+ _02324_ sky130_fd_sc_hd__mux2_1
X_15795_ _08407_ _08408_ vssd1 vssd1 vccd1 vccd1 _08409_ sky130_fd_sc_hd__nor2_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17534_ _09935_ _09938_ _09936_ vssd1 vssd1 vccd1 vccd1 _10071_ sky130_fd_sc_hd__a21bo_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _07358_ _07359_ vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__and2_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_144 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_144/HI o_rgb[2] sky130_fd_sc_hd__conb_1
X_11958_ _04666_ _04667_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__nand2_1
XFILLER_178_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_155 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_155/HI o_rgb[17]
+ sky130_fd_sc_hd__conb_1
XFILLER_83_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17465_ _09848_ _09869_ _10002_ vssd1 vssd1 vccd1 vccd1 _10003_ sky130_fd_sc_hd__a21oi_1
XFILLER_233_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10909_ rbzero.tex_b0\[43\] rbzero.tex_b0\[42\] _03671_ vssd1 vssd1 vccd1 vccd1 _03681_
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14677_ _07312_ vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__clkbuf_1
X_11889_ _04080_ _04599_ _04601_ _04078_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a31o_1
X_19204_ rbzero.spi_registers.new_vshift\[5\] _02775_ vssd1 vssd1 vccd1 vccd1 _02782_
+ sky130_fd_sc_hd__or2_1
XFILLER_242_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16416_ _07890_ _07817_ _07553_ _08893_ vssd1 vssd1 vccd1 vccd1 _09026_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13628_ _05728_ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__buf_2
XFILLER_60_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17396_ _09831_ _09834_ _09830_ vssd1 vssd1 vccd1 vccd1 _09934_ sky130_fd_sc_hd__a21bo_1
XFILLER_193_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19135_ _02727_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__buf_2
X_16347_ _08840_ _08957_ vssd1 vssd1 vccd1 vccd1 _08958_ sky130_fd_sc_hd__xnor2_4
X_13559_ _06236_ _06246_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__or2_1
XFILLER_121_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19066_ _02695_ vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__clkbuf_1
X_16278_ _08274_ _07598_ _08888_ vssd1 vssd1 vccd1 vccd1 _08889_ sky130_fd_sc_hd__or3_1
XFILLER_172_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18017_ _01646_ _01647_ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__nor2_1
XFILLER_86_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15229_ _07842_ vssd1 vssd1 vccd1 vccd1 _07843_ sky130_fd_sc_hd__buf_4
XFILLER_172_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout107 net108 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__buf_2
Xfanout118 net122 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__buf_2
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout129 net140 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_2
XFILLER_214_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19968_ _03119_ vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__clkinv_2
XFILLER_99_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18919_ _02607_ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__clkbuf_4
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19899_ _03112_ vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__clkinv_2
XFILLER_228_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20812_ _00030_ _00828_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20743_ net107 _00759_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20674_ net68 _00690_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21226_ _00275_ _01242_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21157_ _00206_ _01173_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20108_ rbzero.traced_texa\[-10\] rbzero.texV\[-10\] vssd1 vssd1 vccd1 vccd1 _03144_
+ sky130_fd_sc_hd__nor2_1
XFILLER_28_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21088_ _00137_ _01104_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_77_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12930_ _05611_ _05615_ _05618_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__o21a_1
XFILLER_4_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20039_ _03127_ vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__clkinv_2
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _05493_ _05507_ _05478_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__mux2_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _05020_ _07254_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__nor2_1
XFILLER_57_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _04522_ _04525_ _03919_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__mux2_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _08133_ _08142_ vssd1 vssd1 vccd1 vccd1 _08194_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12792_ _05404_ _05445_ _05470_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__a21o_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14531_ rbzero.wall_tracer.stepDistY\[1\] _07206_ _07193_ vssd1 vssd1 vccd1 vccd1
+ _07207_ sky130_fd_sc_hd__mux2_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _04456_ _04457_ _04323_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__mux2_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17250_ _09677_ _09694_ _09692_ vssd1 vssd1 vccd1 vccd1 _09789_ sky130_fd_sc_hd__a21o_1
XFILLER_202_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _07148_ vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11674_ _03958_ _04387_ _04388_ _04389_ _04007_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__o221a_1
XFILLER_202_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16201_ _08810_ _08812_ vssd1 vssd1 vccd1 vccd1 _08813_ sky130_fd_sc_hd__xor2_1
X_13413_ _05671_ _05629_ _05622_ _06101_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__or4_1
XFILLER_70_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17181_ _08787_ _09207_ _08272_ vssd1 vssd1 vccd1 vccd1 _09721_ sky130_fd_sc_hd__a21oi_2
X_10625_ _03532_ vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14393_ _07005_ _07081_ _06990_ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__mux2_1
X_16132_ _08728_ _08743_ vssd1 vssd1 vccd1 vccd1 _08744_ sky130_fd_sc_hd__xor2_1
XFILLER_183_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13344_ _06030_ _06031_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__xor2_1
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10556_ rbzero.tex_r0\[19\] rbzero.tex_r0\[18\] _03490_ vssd1 vssd1 vccd1 vccd1 _03496_
+ sky130_fd_sc_hd__mux2_1
XFILLER_154_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16063_ _08508_ _08511_ _08506_ vssd1 vssd1 vccd1 vccd1 _08676_ sky130_fd_sc_hd__a21bo_1
XFILLER_154_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13275_ _05537_ _05622_ _05886_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__o21ai_1
X_10487_ rbzero.tex_r0\[52\] rbzero.tex_r0\[51\] _03457_ vssd1 vssd1 vccd1 vccd1 _03460_
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15014_ _07518_ _07530_ _07627_ vssd1 vssd1 vccd1 vccd1 _07628_ sky130_fd_sc_hd__a21o_1
X_12226_ _04925_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__buf_4
XFILLER_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12157_ _04853_ _04861_ _04863_ _04860_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__a22o_1
XFILLER_116_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19822_ _03105_ vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__clkinv_2
XFILLER_190_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11108_ rbzero.traced_texVinit\[6\] rbzero.spi_registers.vshift\[3\] vssd1 vssd1
+ vccd1 vccd1 _03827_ sky130_fd_sc_hd__nand2_1
X_16965_ _09369_ _09506_ vssd1 vssd1 vccd1 vccd1 _09507_ sky130_fd_sc_hd__xor2_4
X_12088_ _04775_ _04792_ _04794_ _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__and4_1
X_19753_ rbzero.pov.ready_buffer\[3\] _03069_ _03070_ rbzero.debug_overlay.vplaneY\[-6\]
+ _02832_ vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__o221a_1
XFILLER_46_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15916_ _07902_ _07875_ vssd1 vssd1 vccd1 vccd1 _08530_ sky130_fd_sc_hd__or2b_1
X_11039_ rbzero.otherx\[1\] _03735_ _03746_ rbzero.otherx\[3\] vssd1 vssd1 vccd1 vccd1
+ _03767_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18704_ _02429_ _02430_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__nor2_1
X_19684_ rbzero.pov.ready_buffer\[55\] _02958_ _03007_ _03041_ vssd1 vssd1 vccd1 vccd1
+ _03042_ sky130_fd_sc_hd__a211o_1
XFILLER_237_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16896_ _09436_ _09437_ vssd1 vssd1 vccd1 vccd1 _09438_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18635_ rbzero.map_rom.i_col\[4\] _02367_ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15847_ _07863_ _07865_ _07748_ _07862_ vssd1 vssd1 vccd1 vccd1 _08461_ sky130_fd_sc_hd__a2bb2o_1
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18566_ _02191_ _02291_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__nand2_1
XFILLER_206_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15778_ _08390_ _08391_ vssd1 vssd1 vccd1 vccd1 _08392_ sky130_fd_sc_hd__xnor2_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17517_ _07420_ _07421_ _09389_ vssd1 vssd1 vccd1 vccd1 _10054_ sky130_fd_sc_hd__and3_2
XFILLER_166_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14729_ _07342_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__clkbuf_4
XFILLER_33_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18497_ _02234_ _02235_ _02243_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__o21ai_1
XFILLER_127_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17448_ _09983_ _09984_ _09975_ vssd1 vssd1 vccd1 vccd1 _09986_ sky130_fd_sc_hd__a21oi_1
XFILLER_221_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17379_ _09915_ _09916_ vssd1 vssd1 vccd1 vccd1 _09917_ sky130_fd_sc_hd__or2b_1
XFILLER_159_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19118_ rbzero.spi_registers.new_other\[7\] _02725_ vssd1 vssd1 vccd1 vccd1 _02729_
+ sky130_fd_sc_hd__or2_1
XFILLER_203_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20390_ net135 _00421_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19049_ rbzero.pov.spi_buffer\[71\] rbzero.pov.ready_buffer\[71\] _02607_ vssd1 vssd1
+ vccd1 vccd1 _02686_ sky130_fd_sc_hd__mux2_1
XFILLER_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21011_ net81 _01027_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20726_ net101 _00742_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.vinf sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20657_ net63 _00673_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10410_ _03417_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_149_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11390_ _04101_ _04103_ _04105_ _04106_ _04108_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__o221ai_4
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20588_ net90 _00604_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10341_ rbzero.tex_r1\[54\] rbzero.tex_r1\[55\] _03377_ vssd1 vssd1 vccd1 vccd1 _03381_
+ sky130_fd_sc_hd__mux2_1
XFILLER_164_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13060_ _05567_ _05748_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__nand2_2
X_10272_ rbzero.tex_b1\[23\] rbzero.tex_b1\[24\] _03344_ vssd1 vssd1 vccd1 vccd1 _03345_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12011_ net8 net7 vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__nor2_1
XFILLER_79_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21209_ _00258_ _01225_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16750_ _09275_ vssd1 vssd1 vccd1 vccd1 _09301_ sky130_fd_sc_hd__clkbuf_4
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13962_ _06313_ _06422_ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__nor2_1
XFILLER_47_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15701_ _08188_ _08215_ vssd1 vssd1 vccd1 vccd1 _08315_ sky130_fd_sc_hd__xnor2_2
X_12913_ _05480_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__clkbuf_2
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16681_ rbzero.row_render.texu\[5\] _09260_ _09258_ rbzero.wall_tracer.texu\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__a22o_1
X_13893_ _06578_ _06579_ _06581_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__o21a_1
XFILLER_62_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18420_ rbzero.debug_overlay.vplaneX\[-3\] rbzero.wall_tracer.rayAddendX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__nor2_1
X_15632_ _08231_ _08239_ _08243_ vssd1 vssd1 vccd1 vccd1 _08246_ sky130_fd_sc_hd__or3_1
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _05480_ _05532_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__and2_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _05121_ _02110_ _02111_ _02000_ vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__a31o_1
XFILLER_163_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15563_ _08174_ _08175_ _08176_ vssd1 vssd1 vccd1 vccd1 _08177_ sky130_fd_sc_hd__a21boi_1
XFILLER_15_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _05375_ _05378_ _05395_ _05381_ _05462_ _05463_ vssd1 vssd1 vccd1 vccd1 _05464_
+ sky130_fd_sc_hd__mux4_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17302_ _09577_ _09706_ vssd1 vssd1 vccd1 vccd1 _09841_ sky130_fd_sc_hd__nand2_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14514_ rbzero.wall_tracer.stepDistY\[-3\] _07192_ _07193_ vssd1 vssd1 vccd1 vccd1
+ _07194_ sky130_fd_sc_hd__mux2_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ rbzero.wall_tracer.trackDistY\[-3\] rbzero.wall_tracer.stepDistY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__or2_1
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _03956_ _04429_ _04433_ _04441_ _03985_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__o311a_1
X_15494_ _08073_ _08106_ _08107_ vssd1 vssd1 vccd1 vccd1 _08108_ sky130_fd_sc_hd__a21boi_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17233_ rbzero.wall_tracer.trackDistX\[2\] _09301_ _09765_ _09772_ vssd1 vssd1 vccd1
+ vccd1 _00555_ sky130_fd_sc_hd__o22a_1
XFILLER_202_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14445_ _05538_ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__clkbuf_4
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11657_ _04373_ vssd1 vssd1 vccd1 vccd1 o_rgb[14] sky130_fd_sc_hd__buf_4
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17164_ _07631_ _07760_ vssd1 vssd1 vccd1 vccd1 _09704_ sky130_fd_sc_hd__nor2_1
XFILLER_200_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10608_ _03523_ vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14376_ _06985_ _07032_ _07033_ vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__or3_1
X_11588_ _04303_ _04304_ _03942_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__mux2_1
X_16115_ _08721_ _08726_ vssd1 vssd1 vccd1 vccd1 _08727_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13327_ _05997_ _06014_ _06015_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__a21o_1
XFILLER_122_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17095_ _09514_ _09515_ _09635_ vssd1 vssd1 vccd1 vccd1 _09636_ sky130_fd_sc_hd__and3_1
XFILLER_171_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10539_ rbzero.tex_r0\[27\] rbzero.tex_r0\[26\] _03479_ vssd1 vssd1 vccd1 vccd1 _03487_
+ sky130_fd_sc_hd__mux2_1
X_16046_ _08544_ _08545_ _08546_ _08532_ vssd1 vssd1 vccd1 vccd1 _08659_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_192_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13258_ _05615_ _05939_ _05946_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__a21bo_1
XFILLER_131_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12209_ _04871_ net35 _04911_ _04914_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__a31o_1
XFILLER_83_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13189_ _05842_ _05877_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19805_ _04104_ _04106_ _04113_ _02718_ _03084_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__a41o_1
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17997_ _01777_ _01778_ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__and2_1
XFILLER_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16948_ _09217_ _09218_ vssd1 vssd1 vccd1 vccd1 _09490_ sky130_fd_sc_hd__nor2_1
X_19736_ _03055_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__clkbuf_4
XFILLER_111_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16879_ _09384_ _09179_ _09419_ vssd1 vssd1 vccd1 vccd1 _09421_ sky130_fd_sc_hd__or3_1
X_19667_ rbzero.debug_overlay.playerY\[-2\] _03016_ _03028_ _02978_ vssd1 vssd1 vccd1
+ vccd1 _00982_ sky130_fd_sc_hd__o211a_1
XFILLER_77_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18618_ _03736_ _07491_ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19598_ _02956_ _02974_ _02975_ _02780_ vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__o211a_1
XFILLER_20_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18549_ _02247_ rbzero.debug_overlay.vplaneX\[-2\] vssd1 vssd1 vccd1 vccd1 _02292_
+ sky130_fd_sc_hd__and2_1
XFILLER_212_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20511_ net128 _00527_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20442_ net138 _00473_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_165_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20373_ net118 _00011_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rcp_sel\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_140_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10890_ _03604_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__clkbuf_4
XFILLER_232_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12560_ _05247_ _05248_ _05219_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__mux2_2
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11511_ _03293_ _04228_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__nand2_1
XFILLER_19_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20709_ net84 _00725_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.mosi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12491_ _05178_ _05179_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__nand2_2
XFILLER_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14230_ _06918_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__inv_2
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11442_ _04158_ _04159_ _04014_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__mux2_1
XFILLER_221_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14161_ _06827_ _06849_ vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__nand2_1
X_11373_ _04078_ _04079_ _04077_ _03780_ _04091_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__o221a_1
XFILLER_165_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13112_ _05791_ _05799_ _05800_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__a21o_1
XFILLER_30_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10324_ rbzero.tex_r1\[62\] rbzero.tex_r1\[63\] _03366_ vssd1 vssd1 vccd1 vccd1 _03372_
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14092_ _06751_ _06779_ _06780_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__a21oi_2
XFILLER_193_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17920_ _01599_ _01601_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__nor2_1
XFILLER_180_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13043_ _05725_ _05731_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__xnor2_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ rbzero.tex_b1\[31\] rbzero.tex_b1\[32\] _03333_ vssd1 vssd1 vccd1 vccd1 _03336_
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17851_ _07886_ _08645_ _01632_ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__o21ai_1
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10186_ _03298_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__clkbuf_4
XTAP_6974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16802_ rbzero.wall_tracer.trackDistX\[-3\] rbzero.wall_tracer.stepDistX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _09347_ sky130_fd_sc_hd__nand2_1
XFILLER_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17782_ _01457_ _01467_ _01565_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__a21o_1
XFILLER_226_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14994_ _07508_ _07550_ _07575_ _07542_ vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__o22ai_1
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16733_ _08449_ _08322_ _09285_ vssd1 vssd1 vccd1 vccd1 _09286_ sky130_fd_sc_hd__a21boi_4
X_19521_ rbzero.pov.spi_buffer\[56\] rbzero.pov.spi_buffer\[57\] _02921_ vssd1 vssd1
+ vccd1 vccd1 _02929_ sky130_fd_sc_hd__mux2_1
XFILLER_219_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13945_ _06172_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__buf_2
XFILLER_47_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19452_ rbzero.pov.spi_buffer\[23\] rbzero.pov.spi_buffer\[24\] _02888_ vssd1 vssd1
+ vccd1 vccd1 _02893_ sky130_fd_sc_hd__mux2_1
XFILLER_228_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16664_ rbzero.row_render.size\[1\] _09255_ _07172_ _09259_ vssd1 vssd1 vccd1 vccd1
+ _00499_ sky130_fd_sc_hd__a22o_1
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13876_ _06404_ _06449_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__and2_1
XFILLER_201_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15615_ _08182_ _08181_ vssd1 vssd1 vccd1 vccd1 _08229_ sky130_fd_sc_hd__and2_1
X_18403_ _03729_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__clkbuf_4
X_12827_ _05444_ _05429_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__or2_1
X_19383_ _02861_ vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__clkinv_2
X_16595_ _07826_ _09197_ _09202_ _09203_ vssd1 vssd1 vccd1 vccd1 _09204_ sky130_fd_sc_hd__nor4_1
XFILLER_37_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18334_ _02090_ _02091_ _02089_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__a21boi_1
XFILLER_72_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15546_ _08148_ _08158_ _08159_ vssd1 vssd1 vccd1 vccd1 _08160_ sky130_fd_sc_hd__a21oi_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12758_ _05446_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__buf_4
XFILLER_128_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18265_ _01997_ _02036_ _02037_ _02013_ vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__a31o_1
XFILLER_147_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11709_ _03994_ _04420_ _04424_ _03900_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__a211o_1
XFILLER_230_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15477_ _08081_ _08089_ vssd1 vssd1 vccd1 vccd1 _08091_ sky130_fd_sc_hd__and2b_1
X_12689_ _05251_ _05377_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__xnor2_4
XFILLER_124_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17216_ _09651_ _09755_ vssd1 vssd1 vccd1 vccd1 _09756_ sky130_fd_sc_hd__xnor2_1
XFILLER_204_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14428_ _05577_ _07110_ _07116_ _05602_ vssd1 vssd1 vccd1 vccd1 _07117_ sky130_fd_sc_hd__a211o_1
XFILLER_147_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18196_ _01835_ _01852_ _01975_ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__a21o_1
XFILLER_239_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17147_ _09679_ _09686_ vssd1 vssd1 vccd1 vccd1 _09687_ sky130_fd_sc_hd__and2_1
XFILLER_200_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14359_ _07046_ _07047_ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__nor2_1
XFILLER_116_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17078_ _09601_ _09618_ vssd1 vssd1 vccd1 vccd1 _09619_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16029_ _07824_ _07680_ vssd1 vssd1 vccd1 vccd1 _08642_ sky130_fd_sc_hd__nor2_1
XFILLER_131_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19719_ _02708_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__buf_2
XFILLER_226_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20991_ net90 _01007_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_226_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20425_ net117 _00456_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20356_ _02727_ _03279_ _03280_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__and3_1
XFILLER_101_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20287_ _03257_ vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__clkinv_2
XTAP_6226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11991_ _04694_ _04696_ _04700_ _04667_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__a22o_1
XFILLER_44_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13730_ _05861_ _06389_ _06391_ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__o21bai_1
XFILLER_29_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10942_ _03698_ vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13661_ _06348_ _06349_ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__or2b_1
XFILLER_232_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10873_ _03662_ vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15400_ _08007_ _08013_ vssd1 vssd1 vccd1 vccd1 _08014_ sky130_fd_sc_hd__xor2_2
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ rbzero.wall_tracer.visualWallDist\[10\] vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__clkinv_2
X_16380_ _08429_ _08724_ _08857_ _08854_ vssd1 vssd1 vccd1 vccd1 _08990_ sky130_fd_sc_hd__o31a_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _06237_ _06244_ vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__and2b_1
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15331_ _07474_ _07942_ _07943_ _07944_ vssd1 vssd1 vccd1 vccd1 _07945_ sky130_fd_sc_hd__nand4_1
XFILLER_34_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12543_ _03815_ _05074_ _05090_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__and3_1
XFILLER_129_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18050_ _01728_ _01729_ _01817_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__a21o_1
XFILLER_157_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15262_ _07747_ _07753_ vssd1 vssd1 vccd1 vccd1 _07876_ sky130_fd_sc_hd__nand2_1
X_12474_ _05161_ _05162_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__nor2_2
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17001_ _09540_ _09541_ vssd1 vssd1 vccd1 vccd1 _09542_ sky130_fd_sc_hd__nor2_1
X_14213_ _06898_ _06901_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__and2_1
XFILLER_123_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11425_ _04142_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__buf_2
X_15193_ _07804_ _07806_ vssd1 vssd1 vccd1 vccd1 _07807_ sky130_fd_sc_hd__nor2_1
XFILLER_172_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_7 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14144_ _06825_ _06831_ _06812_ _06813_ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__o211a_1
XFILLER_197_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11356_ _04046_ _04074_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__nor2_1
XFILLER_126_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10307_ rbzero.tex_b1\[6\] rbzero.tex_b1\[7\] _03355_ vssd1 vssd1 vccd1 vccd1 _03363_
+ sky130_fd_sc_hd__mux2_1
X_14075_ _06470_ _06388_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__nor2_1
X_18952_ _02635_ vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11287_ _03900_ _03993_ _04005_ _03954_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__o211a_1
X_17903_ _01596_ _01597_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__or2b_1
X_13026_ _05635_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__buf_2
XFILLER_239_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10238_ rbzero.tex_b1\[39\] rbzero.tex_b1\[40\] _03322_ vssd1 vssd1 vccd1 vccd1 _03327_
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18883_ _02594_ _02595_ _02590_ vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__and3b_1
XTAP_6760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17834_ _01616_ _01617_ _09275_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__o21a_1
XFILLER_239_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17765_ _01452_ _01455_ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__nand2_1
X_14977_ _07501_ vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__buf_2
XFILLER_130_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19504_ rbzero.pov.spi_buffer\[48\] rbzero.pov.spi_buffer\[49\] _02910_ vssd1 vssd1
+ vccd1 vccd1 _02920_ sky130_fd_sc_hd__mux2_1
X_13928_ _06607_ _06616_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__xor2_1
X_16716_ rbzero.wall_tracer.wall\[1\] rbzero.row_render.wall\[1\] _09269_ vssd1 vssd1
+ vccd1 vccd1 _09271_ sky130_fd_sc_hd__mux2_1
XFILLER_130_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17696_ _01478_ _01479_ _10121_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__a21oi_1
XFILLER_207_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16647_ _04220_ _09244_ vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__nor2_1
X_19435_ rbzero.pov.spi_buffer\[15\] rbzero.pov.spi_buffer\[16\] _02877_ vssd1 vssd1
+ vccd1 vccd1 _02884_ sky130_fd_sc_hd__mux2_1
X_13859_ _06465_ _06522_ _06523_ _06532_ vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__a31o_1
XFILLER_165_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16578_ _09047_ _09185_ _09186_ vssd1 vssd1 vccd1 vccd1 _09187_ sky130_fd_sc_hd__o21a_1
X_19366_ _02859_ vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__clkinv_2
XFILLER_222_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18317_ rbzero.wall_tracer.trackDistY\[2\] rbzero.wall_tracer.stepDistY\[2\] vssd1
+ vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__nand2_1
X_15529_ _08134_ _08141_ vssd1 vssd1 vccd1 vccd1 _08143_ sky130_fd_sc_hd__nor2_1
X_19297_ _02740_ _02833_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__or2_1
XFILLER_31_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18248_ _02015_ _02017_ _02016_ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__a21boi_1
XFILLER_198_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18179_ _01957_ _01958_ vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__xnor2_1
XFILLER_175_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20210_ _03228_ _03229_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21190_ _00239_ _01206_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20141_ rbzero.traced_texa\[-4\] rbzero.texV\[-4\] vssd1 vssd1 vccd1 vccd1 _03171_
+ sky130_fd_sc_hd__nor2_1
XFILLER_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20072_ _03130_ vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__clkinv_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20974_ net63 _00990_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11210_ _03928_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__buf_4
X_20408_ net130 _00439_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_135_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12190_ _04883_ _04519_ net37 net36 vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__o211a_1
XFILLER_108_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21388_ net109 _01404_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11141_ _03853_ _03859_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__nor2_2
XTAP_6001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20339_ rbzero.wall_tracer.rayAddendX\[-7\] _03260_ _09267_ _03270_ vssd1 vssd1 vccd1
+ vccd1 _01412_ sky130_fd_sc_hd__a22o_1
XTAP_6012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11072_ _03795_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__buf_4
XFILLER_122_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14900_ _04932_ _07513_ _03793_ vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__o21ai_1
XFILLER_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880_ _08491_ _08492_ _08483_ vssd1 vssd1 vccd1 vccd1 _08494_ sky130_fd_sc_hd__a21o_1
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14831_ _07202_ _07444_ _07206_ vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__a21o_2
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17550_ _10049_ _10050_ _10086_ vssd1 vssd1 vccd1 vccd1 _10087_ sky130_fd_sc_hd__a21o_1
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14762_ _04935_ _07375_ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__nand2_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ net18 net19 _04682_ net20 vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__o22a_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16501_ _08429_ _08852_ _08980_ vssd1 vssd1 vccd1 vccd1 _09110_ sky130_fd_sc_hd__or3_1
XFILLER_229_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13713_ _06400_ _06401_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__xor2_2
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17481_ _10015_ _10017_ vssd1 vssd1 vccd1 vccd1 _10019_ sky130_fd_sc_hd__and2_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10925_ _03689_ vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__clkbuf_1
X_14693_ rbzero.wall_tracer.stepDistX\[1\] _07206_ _07316_ vssd1 vssd1 vccd1 vccd1
+ _07321_ sky130_fd_sc_hd__mux2_1
XFILLER_205_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16432_ _09040_ _09041_ vssd1 vssd1 vccd1 vccd1 _09042_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19220_ _02791_ vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__clkbuf_1
X_13644_ _05722_ _06321_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__and2_1
XFILLER_147_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10856_ _03653_ vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19151_ rbzero.spi_registers.new_leak\[3\] _02745_ vssd1 vssd1 vccd1 vccd1 _02749_
+ sky130_fd_sc_hd__or2_1
X_16363_ _08878_ _08969_ _08971_ vssd1 vssd1 vccd1 vccd1 _08973_ sky130_fd_sc_hd__and3_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _06252_ _06250_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__and2b_1
XFILLER_158_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _03617_ vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18102_ _01630_ _01633_ _01787_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__a21oi_1
XFILLER_197_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _07906_ _07907_ _07927_ vssd1 vssd1 vccd1 vccd1 _07928_ sky130_fd_sc_hd__nand3_1
XFILLER_169_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _05176_ _05214_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__xnor2_2
X_19082_ _02704_ vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__clkbuf_1
X_16294_ _08046_ _08636_ vssd1 vssd1 vccd1 vccd1 _08905_ sky130_fd_sc_hd__nand2_1
XFILLER_184_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18033_ _01700_ vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__inv_2
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15245_ _07469_ _07858_ _07750_ _07749_ vssd1 vssd1 vccd1 vccd1 _07859_ sky130_fd_sc_hd__o31ai_2
X_12457_ rbzero.debug_overlay.facingX\[-1\] rbzero.wall_tracer.rayAddendX\[7\] _05144_
+ _05145_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__a31o_1
X_11408_ _04122_ _04125_ _03923_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__mux2_1
X_15176_ _07510_ vssd1 vssd1 vccd1 vccd1 _07790_ sky130_fd_sc_hd__buf_2
XFILLER_158_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12388_ _05034_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__inv_2
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14127_ _06815_ _06801_ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__xor2_1
XFILLER_99_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11339_ _04056_ gpout0.hpos\[1\] gpout0.hpos\[0\] _04057_ vssd1 vssd1 vccd1 vccd1
+ _04058_ sky130_fd_sc_hd__o211a_1
XFILLER_99_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19984_ _03121_ vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__clkinv_2
XFILLER_207_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14058_ _06698_ _06742_ _06746_ vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__a21boi_1
X_18935_ _02626_ vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13009_ _05666_ _05697_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__xor2_1
XFILLER_136_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18866_ rbzero.spi_registers.spi_cmd\[2\] vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__inv_2
XTAP_6590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17817_ _01448_ _01487_ _01600_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__a21oi_1
XFILLER_227_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18797_ _02505_ _02513_ _02517_ vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__nand3_1
XFILLER_48_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17748_ _08135_ _09115_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__nor2_1
XFILLER_236_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17679_ _01462_ _01463_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19418_ rbzero.pov.spi_buffer\[7\] rbzero.pov.spi_buffer\[8\] _02866_ vssd1 vssd1
+ vccd1 vccd1 _02875_ sky130_fd_sc_hd__mux2_1
X_20690_ net70 _00706_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[70\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19349_ _02855_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__buf_4
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21311_ net112 _01327_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21242_ _00291_ _01258_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21173_ _00222_ _01189_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20124_ _03093_ _03156_ _03157_ _03137_ rbzero.texV\[-8\] vssd1 vssd1 vccd1 vccd1
+ _01310_ sky130_fd_sc_hd__a32o_1
XFILLER_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20055_ _03128_ vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__clkinv_2
XFILLER_98_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ net70 _00973_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ rbzero.tex_g1\[9\] rbzero.tex_g1\[10\] _03574_ vssd1 vssd1 vccd1 vccd1 _03577_
+ sky130_fd_sc_hd__mux2_1
XFILLER_187_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _04323_ _04403_ _04404_ _04405_ _03972_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__o221a_1
XFILLER_198_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20888_ net62 _00904_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10641_ _03540_ vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13360_ _06047_ _06048_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__or2b_1
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10572_ _03504_ vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12311_ rbzero.wall_tracer.trackDistX\[7\] _04999_ rbzero.wall_tracer.trackDistX\[6\]
+ _05004_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__o22a_1
XFILLER_158_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13291_ _05978_ _05979_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__and2_1
XFILLER_108_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15030_ rbzero.debug_overlay.playerX\[-9\] rbzero.wall_tracer.state\[6\] _07643_
+ vssd1 vssd1 vccd1 vccd1 _07644_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12242_ _04935_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__buf_4
XFILLER_68_1322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12173_ net36 _04878_ _04873_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__o21ba_1
XFILLER_194_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11124_ rbzero.traced_texVinit\[4\] rbzero.spi_registers.vshift\[1\] vssd1 vssd1
+ vccd1 vccd1 _03843_ sky130_fd_sc_hd__or2_1
XFILLER_96_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16981_ _09520_ _09521_ vssd1 vssd1 vccd1 vccd1 _09522_ sky130_fd_sc_hd__or2_1
XFILLER_150_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18720_ _02442_ _02443_ _02444_ _02445_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__nand4_2
X_15932_ _08544_ _08545_ vssd1 vssd1 vccd1 vccd1 _08546_ sky130_fd_sc_hd__xor2_1
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11055_ gpout0.hpos\[3\] gpout0.hpos\[4\] vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__and2_1
XFILLER_114_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15863_ _04933_ _08474_ _08476_ _07822_ vssd1 vssd1 vccd1 vccd1 _08477_ sky130_fd_sc_hd__a31o_1
XTAP_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18651_ _02371_ _02372_ _02382_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__or3_1
XFILLER_188_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ _10047_ _10138_ vssd1 vssd1 vccd1 vccd1 _10139_ sky130_fd_sc_hd__xnor2_1
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14814_ _07427_ rbzero.debug_overlay.playerY\[-8\] _05113_ vssd1 vssd1 vccd1 vccd1
+ _07428_ sky130_fd_sc_hd__mux2_1
XFILLER_224_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15794_ _08380_ _08375_ _08379_ vssd1 vssd1 vccd1 vccd1 _08408_ sky130_fd_sc_hd__a21oi_1
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18582_ _02318_ _02319_ _03818_ _02322_ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_236_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17533_ _10068_ _10069_ vssd1 vssd1 vccd1 vccd1 _10070_ sky130_fd_sc_hd__and2_1
X_14745_ rbzero.debug_overlay.playerY\[-6\] _07357_ vssd1 vssd1 vccd1 vccd1 _07359_
+ sky130_fd_sc_hd__nand2_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ net20 net19 vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__nor2_1
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_145 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_145/HI o_rgb[3] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_156 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_156/HI o_rgb[18]
+ sky130_fd_sc_hd__conb_1
XFILLER_229_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17464_ _09866_ _09868_ vssd1 vssd1 vccd1 vccd1 _10002_ sky130_fd_sc_hd__and2_1
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10908_ _03680_ vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__clkbuf_1
XFILLER_205_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14676_ rbzero.wall_tracer.stepDistX\[-7\] _07172_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _07312_ sky130_fd_sc_hd__mux2_1
X_11888_ _04600_ _04591_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__or2b_1
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16415_ _07890_ _07800_ _07685_ _07817_ vssd1 vssd1 vccd1 vccd1 _09025_ sky130_fd_sc_hd__or4_1
X_19203_ rbzero.spi_registers.vshift\[4\] _02774_ _02781_ _02780_ vssd1 vssd1 vccd1
+ vccd1 _00765_ sky130_fd_sc_hd__o211a_1
X_13627_ _06309_ _06315_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__nor2_1
XFILLER_177_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17395_ _09811_ _09813_ _09810_ vssd1 vssd1 vccd1 vccd1 _09933_ sky130_fd_sc_hd__a21bo_1
XFILLER_158_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10839_ _03644_ vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16346_ _08955_ _08956_ vssd1 vssd1 vccd1 vccd1 _08957_ sky130_fd_sc_hd__and2_2
XFILLER_158_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19134_ rbzero.spi_registers.new_other\[4\] _02725_ vssd1 vssd1 vccd1 vccd1 _02737_
+ sky130_fd_sc_hd__or2_1
XFILLER_203_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13558_ _06236_ _06246_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__nand2_1
XFILLER_242_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12509_ _05071_ _05072_ _03815_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__and3b_1
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19065_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.spi_buffer\[3\]
+ _02690_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__mux2_1
X_16277_ _08886_ _08887_ vssd1 vssd1 vccd1 vccd1 _08888_ sky130_fd_sc_hd__nand2_1
X_13489_ _05877_ _05842_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__and2b_1
XFILLER_51_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18016_ _01756_ _01797_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15228_ _07841_ vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__buf_2
XFILLER_12_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15159_ _07757_ _07772_ vssd1 vssd1 vccd1 vccd1 _07773_ sky130_fd_sc_hd__xor2_1
XFILLER_173_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout108 net141 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__buf_2
XFILLER_99_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout119 net122 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__buf_2
X_19967_ _03119_ vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__clkinv_2
XFILLER_141_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18918_ _02617_ vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19898_ _03112_ vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__clkinv_2
XFILLER_214_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18849_ _02563_ _02564_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__or2_1
XFILLER_216_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20811_ _00029_ _00827_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20742_ net106 _00758_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20673_ net68 _00689_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21225_ _00274_ _01241_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21156_ _00205_ _01172_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20107_ _03139_ _03140_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__and2_1
XFILLER_24_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21087_ _00136_ _01103_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20038_ _03127_ vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__clkinv_2
XFILLER_59_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ _05405_ _05548_ _05504_ _05406_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__o2bb2a_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _04523_ _04524_ _03928_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__mux2_1
XFILLER_233_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _05416_ _05360_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__nand2_2
XFILLER_61_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _07099_ _07204_ _07205_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__nand3_4
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ rbzero.tex_b0\[51\] rbzero.tex_b0\[50\] _04013_ vssd1 vssd1 vccd1 vccd1 _04457_
+ sky130_fd_sc_hd__mux2_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ rbzero.wall_tracer.stepDistY\[-10\] _07147_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _07148_ sky130_fd_sc_hd__mux2_1
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ rbzero.tex_g1\[23\] _03964_ _03965_ _03997_ vssd1 vssd1 vccd1 vccd1 _04389_
+ sky130_fd_sc_hd__a31o_1
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16200_ _08614_ _08655_ _08811_ vssd1 vssd1 vccd1 vccd1 _08812_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13412_ _05631_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__clkbuf_4
X_17180_ _08771_ _09055_ vssd1 vssd1 vccd1 vccd1 _09720_ sky130_fd_sc_hd__and2_1
X_10624_ rbzero.tex_g1\[50\] rbzero.tex_g1\[51\] _03530_ vssd1 vssd1 vccd1 vccd1 _03532_
+ sky130_fd_sc_hd__mux2_1
X_14392_ _07023_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__clkinv_2
XFILLER_126_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16131_ _08741_ _08742_ vssd1 vssd1 vccd1 vccd1 _08743_ sky130_fd_sc_hd__nor2_1
XFILLER_155_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13343_ _05671_ _05746_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__nor2_1
XFILLER_167_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10555_ _03495_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16062_ _08673_ _08674_ vssd1 vssd1 vccd1 vccd1 _08675_ sky130_fd_sc_hd__xor2_1
XFILLER_143_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13274_ _05537_ _05622_ _05886_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__or3_1
X_10486_ _03459_ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15013_ _07623_ _07626_ vssd1 vssd1 vccd1 vccd1 _07627_ sky130_fd_sc_hd__or2_1
X_12225_ _04924_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__clkbuf_4
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19821_ _03105_ vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__clkinv_2
XFILLER_68_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12156_ net51 _04848_ _04849_ net53 _04862_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__a221o_1
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11107_ _03825_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__clkinv_2
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19752_ rbzero.pov.ready_buffer\[2\] _03069_ _03070_ rbzero.debug_overlay.vplaneY\[-7\]
+ _02832_ vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__o221a_1
XFILLER_231_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16964_ _09504_ _09505_ vssd1 vssd1 vccd1 vccd1 _09506_ sky130_fd_sc_hd__nor2_2
X_12087_ net24 net25 _04793_ net26 vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__o22a_1
XFILLER_46_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18703_ rbzero.debug_overlay.vplaneY\[0\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__and2_1
X_15915_ _08527_ _08528_ vssd1 vssd1 vccd1 vccd1 _08529_ sky130_fd_sc_hd__xor2_1
X_11038_ rbzero.othery\[4\] vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__inv_2
XFILLER_231_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19683_ _03039_ _03040_ _02835_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__a21oi_1
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16895_ _07805_ _07817_ vssd1 vssd1 vccd1 vccd1 _09437_ sky130_fd_sc_hd__or2_1
XFILLER_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18634_ _07491_ _02356_ _02366_ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__o21ai_1
X_15846_ _07961_ _08034_ vssd1 vssd1 vccd1 vccd1 _08460_ sky130_fd_sc_hd__nor2_1
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18565_ _02305_ _02306_ _02291_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__o21bai_1
X_15777_ _07792_ _07843_ vssd1 vssd1 vccd1 vccd1 _08391_ sky130_fd_sc_hd__nor2_1
X_12989_ _05621_ _05631_ _05641_ _05645_ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__a2bb2o_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17516_ _10051_ _10052_ vssd1 vssd1 vccd1 vccd1 _10053_ sky130_fd_sc_hd__nand2_1
X_14728_ _07341_ vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__buf_2
XFILLER_127_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18496_ _02241_ _02242_ _03811_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__o21a_1
XFILLER_33_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17447_ _09975_ _09983_ _09984_ vssd1 vssd1 vccd1 vccd1 _09985_ sky130_fd_sc_hd__and3_1
X_14659_ rbzero.wall_tracer.visualWallDist\[9\] _07252_ vssd1 vssd1 vccd1 vccd1 _07303_
+ sky130_fd_sc_hd__or2_1
XFILLER_177_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17378_ _08890_ _08596_ _08850_ _08978_ vssd1 vssd1 vccd1 vccd1 _09916_ sky130_fd_sc_hd__or4_1
XFILLER_193_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19117_ rbzero.otherx\[0\] _02723_ _02726_ _02728_ vssd1 vssd1 vccd1 vccd1 _00732_
+ sky130_fd_sc_hd__o211a_1
X_16329_ _08937_ _08939_ vssd1 vssd1 vccd1 vccd1 _08940_ sky130_fd_sc_hd__xor2_1
XFILLER_174_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19048_ _02685_ vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21010_ net80 _01026_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_86_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20725_ net101 _00741_ vssd1 vssd1 vccd1 vccd1 rbzero.othery\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20656_ net63 _00672_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_221_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20587_ net90 _00603_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_221_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10340_ _03380_ vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10271_ _03299_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__clkbuf_4
XFILLER_105_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12010_ net5 net6 vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__nor2_1
XFILLER_156_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21208_ _00257_ _01224_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21139_ _00188_ _01155_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13961_ _06266_ _06483_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__or2_1
XFILLER_4_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15700_ _08283_ _08312_ _08313_ vssd1 vssd1 vccd1 vccd1 _08314_ sky130_fd_sc_hd__a21oi_1
X_12912_ _05501_ _05560_ _05600_ _05405_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__o211a_1
XFILLER_150_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16680_ rbzero.row_render.texu\[4\] _09260_ _09258_ rbzero.wall_tracer.texu\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__a22o_1
XFILLER_219_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13892_ _05861_ _06172_ _06580_ vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__or3_1
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12843_ _05530_ _05473_ _05531_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__mux2_1
X_15631_ _08191_ _08212_ vssd1 vssd1 vccd1 vccd1 _08245_ sky130_fd_sc_hd__xnor2_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18350_ _02107_ _02108_ _02109_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__o21ai_1
X_15562_ _07435_ _08086_ _07484_ _07970_ vssd1 vssd1 vccd1 vccd1 _08176_ sky130_fd_sc_hd__or4_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12774_ _05448_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__clkbuf_4
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _09838_ _09839_ vssd1 vssd1 vccd1 vccd1 _09840_ sky130_fd_sc_hd__xor2_1
XFILLER_202_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14513_ _04925_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__clkbuf_4
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11725_ _04007_ _04436_ _04440_ _03899_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__a211o_1
X_18281_ rbzero.wall_tracer.trackDistY\[-4\] _02039_ _02051_ _09338_ vssd1 vssd1 vccd1
+ vccd1 _00573_ sky130_fd_sc_hd__o22a_1
XFILLER_163_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15493_ _08074_ _08105_ vssd1 vssd1 vccd1 vccd1 _08107_ sky130_fd_sc_hd__or2b_1
XFILLER_30_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17232_ _09303_ _09770_ _09771_ _09282_ vssd1 vssd1 vccd1 vccd1 _09772_ sky130_fd_sc_hd__a31o_1
X_14444_ _07130_ _07046_ _07131_ _07115_ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__a22o_1
XFILLER_175_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11656_ _03826_ _04372_ _04117_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__o21ba_1
XFILLER_202_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout90 net92 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_2
XFILLER_204_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17163_ _09701_ _09702_ vssd1 vssd1 vccd1 vccd1 _09703_ sky130_fd_sc_hd__and2b_1
X_10607_ rbzero.tex_g1\[58\] rbzero.tex_g1\[59\] _03519_ vssd1 vssd1 vccd1 vccd1 _03523_
+ sky130_fd_sc_hd__mux2_1
X_14375_ _06981_ _06980_ _07030_ _06987_ vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__a211o_1
XFILLER_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11587_ rbzero.tex_g0\[17\] rbzero.tex_g0\[16\] _04119_ vssd1 vssd1 vccd1 vccd1 _04304_
+ sky130_fd_sc_hd__mux2_1
XFILLER_200_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16114_ _07625_ _08725_ vssd1 vssd1 vccd1 vccd1 _08726_ sky130_fd_sc_hd__nor2_1
XFILLER_196_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13326_ _05999_ _06013_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__nor2_1
X_17094_ _09516_ _09634_ vssd1 vssd1 vccd1 vccd1 _09635_ sky130_fd_sc_hd__xor2_1
X_10538_ _03486_ vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16045_ _08656_ _08657_ vssd1 vssd1 vccd1 vccd1 _08658_ sky130_fd_sc_hd__xor2_1
XFILLER_170_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13257_ _05940_ _05945_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__or2b_1
X_10469_ _03450_ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12208_ _04885_ _04913_ net38 vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__a21o_1
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13188_ _05874_ _05876_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__xor2_1
XFILLER_111_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19804_ gpout0.vpos\[8\] _03099_ _03102_ _03031_ vssd1 vssd1 vccd1 vccd1 _01045_
+ sky130_fd_sc_hd__o211a_1
X_12139_ net30 net31 _04844_ net32 vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__o22a_1
X_17996_ _01766_ _01776_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__or2_1
XFILLER_111_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19735_ rbzero.pov.ready_buffer\[31\] _03067_ _03068_ rbzero.debug_overlay.facingY\[0\]
+ _03066_ vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__a221o_1
X_16947_ _09446_ _09488_ vssd1 vssd1 vccd1 vccd1 _09489_ sky130_fd_sc_hd__xnor2_1
XFILLER_211_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19666_ _07543_ _02836_ _03016_ _03027_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__o211ai_1
X_16878_ _09384_ _09179_ _09419_ vssd1 vssd1 vccd1 vccd1 _09420_ sky130_fd_sc_hd__o21ai_1
XFILLER_42_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18617_ _02352_ vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15829_ _08351_ _08352_ vssd1 vssd1 vccd1 vccd1 _08443_ sky130_fd_sc_hd__xor2_1
XFILLER_20_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19597_ _07537_ _02960_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__nand2_1
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18548_ _02274_ rbzero.debug_overlay.vplaneX\[-2\] vssd1 vssd1 vccd1 vccd1 _02291_
+ sky130_fd_sc_hd__nor2_1
XFILLER_240_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18479_ _02212_ _02215_ _02225_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__nand3_1
XFILLER_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20510_ net132 _00526_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20441_ net138 _00472_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20372_ net97 _00405_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.i_row\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11510_ _04205_ _04204_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__and2b_1
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20708_ net99 _00724_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12490_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[9\] vssd1
+ vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__nand2_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11441_ rbzero.tex_r1\[17\] rbzero.tex_r1\[16\] _04148_ vssd1 vssd1 vccd1 vccd1 _04159_
+ sky130_fd_sc_hd__mux2_1
X_20639_ net56 _00655_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14160_ _06743_ _06804_ vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__or2_1
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11372_ _04080_ _04082_ _04079_ gpout0.hpos\[4\] _04090_ vssd1 vssd1 vccd1 vccd1
+ _04091_ sky130_fd_sc_hd__a221o_1
XFILLER_192_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13111_ _05794_ _05798_ _05792_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__o21a_1
XFILLER_137_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10323_ _03371_ vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__clkbuf_1
X_14091_ _06752_ _06778_ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__and2b_1
XFILLER_125_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13042_ _05715_ _05726_ _05729_ _05730_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__o31a_1
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10254_ _03335_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17850_ _07886_ _08645_ _01632_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__or3_1
XFILLER_182_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10185_ _03289_ _03291_ _03292_ _03297_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__and4_2
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16801_ rbzero.wall_tracer.trackDistX\[-3\] rbzero.wall_tracer.stepDistX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _09346_ sky130_fd_sc_hd__or2_1
XTAP_6997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17781_ _01464_ _01466_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__nor2_1
XFILLER_78_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14993_ _07606_ vssd1 vssd1 vccd1 vccd1 _07607_ sky130_fd_sc_hd__inv_2
XFILLER_120_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19520_ _02928_ vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16732_ _08449_ _08322_ _04940_ vssd1 vssd1 vccd1 vccd1 _09285_ sky130_fd_sc_hd__o21a_1
XFILLER_247_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13944_ _06602_ _06620_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19451_ _02892_ vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__clkbuf_1
X_13875_ _06456_ _06503_ vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__nor2_1
XFILLER_189_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16663_ rbzero.row_render.size\[0\] _09255_ _07165_ _09259_ vssd1 vssd1 vccd1 vccd1
+ _00498_ sky130_fd_sc_hd__a22o_1
XFILLER_235_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18402_ _02145_ _02155_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15614_ _07697_ _07579_ _08224_ _08226_ _08227_ vssd1 vssd1 vccd1 vccd1 _08228_ sky130_fd_sc_hd__a32oi_4
X_12826_ _05444_ _05463_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__nand2_1
XFILLER_62_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19382_ _02855_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__buf_4
X_16594_ _07843_ _09051_ _09200_ _08398_ vssd1 vssd1 vccd1 vccd1 _09203_ sky130_fd_sc_hd__o22a_1
XFILLER_188_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18333_ rbzero.wall_tracer.trackDistY\[4\] rbzero.wall_tracer.stepDistY\[4\] vssd1
+ vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__and2_1
XFILLER_203_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12757_ _05404_ _05445_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__and2_1
X_15545_ _08116_ _08147_ vssd1 vssd1 vccd1 vccd1 _08159_ sky130_fd_sc_hd__nor2_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11708_ _04421_ _04422_ _04423_ _03958_ _04007_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__o221a_1
XFILLER_163_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15476_ _08081_ _08089_ vssd1 vssd1 vccd1 vccd1 _08090_ sky130_fd_sc_hd__xnor2_1
X_18264_ _02033_ _02034_ _02035_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__o21ai_1
X_12688_ _05253_ _05255_ _05305_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__o21ai_2
XFILLER_129_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17215_ _09752_ _09754_ vssd1 vssd1 vccd1 vccd1 _09755_ sky130_fd_sc_hd__xor2_1
X_14427_ _07107_ _07113_ _07114_ _07115_ _05577_ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__a221oi_1
XFILLER_175_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ rbzero.tex_g0\[45\] rbzero.tex_g0\[44\] _04000_ vssd1 vssd1 vccd1 vccd1 _04356_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18195_ _01853_ _01888_ vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__and2b_1
XFILLER_128_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17146_ _09683_ _09685_ vssd1 vssd1 vccd1 vccd1 _09686_ sky130_fd_sc_hd__xnor2_1
X_14358_ _05593_ _07010_ vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__nor2_1
XFILLER_239_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13309_ _05965_ _05966_ _05962_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__a21oi_1
X_17077_ _09615_ _09617_ vssd1 vssd1 vccd1 vccd1 _09618_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14289_ _06370_ _06977_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__nand2_1
XFILLER_171_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16028_ _07696_ _08640_ _07835_ vssd1 vssd1 vccd1 vccd1 _08641_ sky130_fd_sc_hd__a21oi_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17979_ _07670_ _08851_ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__or2_1
XFILLER_66_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19718_ rbzero.pov.ready_buffer\[39\] _03061_ _03063_ rbzero.debug_overlay.facingX\[-3\]
+ _03064_ vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__a221o_1
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20990_ net66 _01006_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19649_ _03012_ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__buf_2
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20424_ net124 _00455_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20355_ gpout2.clk_div\[0\] gpout2.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__or2_1
XFILLER_162_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20286_ _03257_ vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__clkinv_2
XFILLER_66_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11990_ net51 _04697_ _04698_ net53 _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__a221o_1
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10941_ rbzero.tex_b0\[28\] rbzero.tex_b0\[27\] _03693_ vssd1 vssd1 vccd1 vccd1 _03698_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13660_ _06329_ _06337_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10872_ rbzero.tex_b0\[61\] rbzero.tex_b0\[60\] _03660_ vssd1 vssd1 vccd1 vccd1 _03662_
+ sky130_fd_sc_hd__mux2_1
XFILLER_232_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12611_ _05292_ _05299_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__xnor2_1
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13591_ _06247_ _06279_ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__xnor2_1
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15330_ _07468_ _07469_ _07456_ _07473_ vssd1 vssd1 vccd1 vccd1 _07944_ sky130_fd_sc_hd__a2bb2o_1
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ rbzero.wall_tracer.visualWallDist\[-5\] _05189_ rbzero.wall_tracer.rcp_sel\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__a21o_1
XFILLER_160_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15261_ _07798_ _07808_ _07807_ vssd1 vssd1 vccd1 vccd1 _07875_ sky130_fd_sc_hd__a21o_1
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12473_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] vssd1
+ vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__nor2_1
X_17000_ _08510_ _08724_ _09394_ _09392_ vssd1 vssd1 vccd1 vccd1 _09541_ sky130_fd_sc_hd__o31a_1
XFILLER_200_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14212_ _06899_ _06900_ vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__nand2_1
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11424_ _03938_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__clkbuf_4
XFILLER_201_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15192_ _07556_ _07805_ _07575_ _07551_ vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__o31a_1
XFILLER_137_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_8 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ _06812_ _06813_ _06825_ _06831_ vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__a211o_1
X_11355_ rbzero.row_render.size\[6\] _04045_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__nor2_1
XFILLER_10_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10306_ _03362_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__clkbuf_1
X_14074_ _06762_ _06720_ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__xnor2_1
XFILLER_180_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18951_ rbzero.pov.spi_buffer\[24\] rbzero.pov.ready_buffer\[24\] _02629_ vssd1 vssd1
+ vccd1 vccd1 _02635_ sky130_fd_sc_hd__mux2_1
XFILLER_193_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11286_ _03994_ _03998_ _04004_ _03956_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__a211o_1
XFILLER_180_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17902_ _01648_ _01684_ vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__xnor2_1
X_13025_ _05703_ _05704_ _05625_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__a21o_1
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10237_ _03326_ vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__clkbuf_1
X_18882_ rbzero.spi_registers.spi_counter\[1\] rbzero.spi_registers.spi_counter\[0\]
+ _02576_ rbzero.spi_registers.spi_counter\[2\] vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a31o_1
XTAP_6750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17833_ _01613_ _01614_ _01615_ _09351_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__a31o_1
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17764_ _01432_ _01435_ _01433_ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__a21bo_1
X_14976_ _07588_ _07589_ vssd1 vssd1 vccd1 vccd1 _07590_ sky130_fd_sc_hd__nand2_1
XFILLER_212_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19503_ _02919_ vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16715_ _09270_ vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13927_ _06609_ _06614_ _06615_ vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__a21oi_1
X_17695_ _10121_ _01478_ _01479_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__and3_1
XFILLER_75_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19434_ _02883_ vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__clkbuf_1
XFILLER_228_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16646_ _04196_ _09244_ vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__nor2_1
X_13858_ _06538_ _06546_ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__nor2_1
XFILLER_211_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12809_ _05495_ _05496_ _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__mux2_1
X_19365_ _02859_ vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__clkinv_2
XFILLER_76_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16577_ _08398_ _09048_ _09051_ vssd1 vssd1 vccd1 vccd1 _09186_ sky130_fd_sc_hd__or3_1
XFILLER_16_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13789_ _06424_ _06427_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18316_ rbzero.wall_tracer.trackDistY\[1\] _02039_ _02081_ _09641_ vssd1 vssd1 vccd1
+ vccd1 _00578_ sky130_fd_sc_hd__o22a_1
XFILLER_176_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15528_ _08134_ _08141_ vssd1 vssd1 vccd1 vccd1 _08142_ sky130_fd_sc_hd__xor2_1
XFILLER_124_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19296_ net40 net39 vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__nor2_4
XFILLER_203_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18247_ rbzero.wall_tracer.trackDistY\[-8\] rbzero.wall_tracer.stepDistY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__and2_1
X_15459_ _07992_ _08072_ vssd1 vssd1 vccd1 vccd1 _08073_ sky130_fd_sc_hd__nor2_1
XFILLER_129_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18178_ _09955_ _08725_ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__nor2_1
XFILLER_141_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17129_ _09022_ _08890_ _08718_ rbzero.wall_tracer.visualWallDist\[7\] vssd1 vssd1
+ vccd1 vccd1 _09669_ sky130_fd_sc_hd__or4b_1
XFILLER_190_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20140_ rbzero.texV\[-5\] _02989_ _03142_ _03170_ vssd1 vssd1 vccd1 vccd1 _01313_
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20071_ _03130_ vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__clkinv_2
XFILLER_174_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20973_ net91 _00989_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_226_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20407_ net128 _00438_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_120_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21387_ net109 _01403_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_218_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11140_ _03855_ _03858_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__or2_2
XFILLER_190_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20338_ _02151_ _03269_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__xnor2_1
XTAP_6002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11071_ _03794_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__buf_4
XFILLER_62_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20269_ _03255_ vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__clkinv_2
XTAP_5312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14830_ _07099_ _07195_ _07198_ vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__nand3_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14761_ _07340_ _07367_ _07374_ vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__mux2_1
X_11973_ net18 net19 _04682_ net20 vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__a22oi_1
XFILLER_229_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16500_ _09012_ _08975_ vssd1 vssd1 vccd1 vccd1 _09109_ sky130_fd_sc_hd__or2b_1
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _06363_ _06361_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__xnor2_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10924_ rbzero.tex_b0\[36\] rbzero.tex_b0\[35\] _03682_ vssd1 vssd1 vccd1 vccd1 _03689_
+ sky130_fd_sc_hd__mux2_1
XFILLER_244_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17480_ _10015_ _10017_ vssd1 vssd1 vccd1 vccd1 _10018_ sky130_fd_sc_hd__nor2_1
XFILLER_186_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14692_ _07320_ vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__clkbuf_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16431_ _07751_ _07834_ vssd1 vssd1 vccd1 vccd1 _09041_ sky130_fd_sc_hd__nor2_1
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13643_ _05861_ _06331_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__nor2_1
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10855_ rbzero.tex_g0\[5\] rbzero.tex_g0\[4\] _03649_ vssd1 vssd1 vccd1 vccd1 _03653_
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19150_ rbzero.floor_leak\[2\] _02744_ _02748_ _02738_ vssd1 vssd1 vccd1 vccd1 _00745_
+ sky130_fd_sc_hd__o211a_1
X_16362_ _08878_ _08969_ _08971_ vssd1 vssd1 vccd1 vccd1 _08972_ sky130_fd_sc_hd__a21oi_2
X_13574_ _06253_ _06228_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__and2b_1
XFILLER_34_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10786_ rbzero.tex_g0\[38\] rbzero.tex_g0\[37\] _03616_ vssd1 vssd1 vccd1 vccd1 _03617_
+ sky130_fd_sc_hd__mux2_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18101_ _01872_ _01881_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15313_ _07637_ _07926_ vssd1 vssd1 vccd1 vccd1 _07927_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12525_ _05168_ _05171_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__or2_1
X_16293_ _08618_ _08772_ _08773_ _08775_ vssd1 vssd1 vccd1 vccd1 _08904_ sky130_fd_sc_hd__a2bb2o_1
X_19081_ rbzero.spi_registers.mosi rbzero.spi_registers.spi_cmd\[0\] _02703_ vssd1
+ vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__mux2_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18032_ _01812_ _01813_ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15244_ _07751_ vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__clkbuf_4
XFILLER_185_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12456_ rbzero.debug_overlay.facingX\[0\] rbzero.wall_tracer.rayAddendX\[8\] vssd1
+ vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__and2_1
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11407_ _04123_ _04124_ _03942_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__mux2_1
X_15175_ _07505_ _07506_ vssd1 vssd1 vccd1 vccd1 _07789_ sky130_fd_sc_hd__and2_1
XFILLER_158_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12387_ _05063_ _05079_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__xnor2_2
XFILLER_126_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14126_ _06137_ _06423_ _06510_ _06800_ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__o31a_1
XFILLER_126_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11338_ rbzero.row_render.size\[0\] vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__inv_2
XFILLER_99_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19983_ _03121_ vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__clkinv_2
XFILLER_45_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14057_ _06266_ _06172_ _06745_ vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__or3b_1
XFILLER_49_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18934_ rbzero.pov.spi_buffer\[16\] rbzero.pov.ready_buffer\[16\] _02618_ vssd1 vssd1
+ vccd1 vccd1 _02626_ sky130_fd_sc_hd__mux2_1
XFILLER_140_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11269_ rbzero.tex_r0\[17\] rbzero.tex_r0\[16\] _03974_ vssd1 vssd1 vccd1 vccd1 _03988_
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13008_ _05687_ _05695_ _05696_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__a21o_1
XFILLER_80_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18865_ rbzero.spi_registers.spi_counter\[3\] _02579_ rbzero.spi_registers.spi_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__mux2_1
XTAP_6580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17816_ _01485_ _01486_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__nor2_1
XFILLER_227_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18796_ _02472_ rbzero.wall_tracer.rayAddendY\[6\] vssd1 vssd1 vccd1 vccd1 _02517_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_223_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17747_ _01528_ _01529_ _01530_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__a21o_1
XFILLER_130_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14959_ _04927_ rbzero.wall_tracer.stepDistX\[-8\] vssd1 vssd1 vccd1 vccd1 _07573_
+ sky130_fd_sc_hd__nor2_2
XFILLER_48_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17678_ _09968_ _09197_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__nor2_1
XFILLER_74_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19417_ _02874_ vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__clkbuf_1
X_16629_ rbzero.debug_overlay.playerY\[-1\] rbzero.debug_overlay.playerX\[-1\] _07343_
+ vssd1 vssd1 vccd1 vccd1 _09238_ sky130_fd_sc_hd__mux2_1
XFILLER_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19348_ _02857_ vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__clkinv_2
XFILLER_17_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19279_ rbzero.spi_registers.got_new_other _02742_ _02740_ _02813_ vssd1 vssd1 vccd1
+ vccd1 _00799_ sky130_fd_sc_hd__a31o_1
XFILLER_241_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21310_ net112 _01326_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21241_ _00290_ _01257_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21172_ _00221_ _01188_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20123_ _03153_ _03154_ _03155_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__or3_1
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20054_ _03128_ vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__clkinv_2
XFILLER_100_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20956_ net91 _00972_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20887_ net62 _00903_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_241_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10640_ rbzero.tex_g1\[42\] rbzero.tex_g1\[43\] _03530_ vssd1 vssd1 vccd1 vccd1 _03540_
+ sky130_fd_sc_hd__mux2_1
XFILLER_146_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10571_ rbzero.tex_r0\[12\] rbzero.tex_r0\[11\] _03501_ vssd1 vssd1 vccd1 vccd1 _03504_
+ sky130_fd_sc_hd__mux2_1
XFILLER_220_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12310_ rbzero.wall_tracer.trackDistY\[6\] vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__inv_2
XFILLER_166_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13290_ _05933_ _05932_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12241_ rbzero.wall_tracer.state\[6\] vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__buf_2
XFILLER_108_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12172_ _03294_ _03295_ gpout0.vpos\[8\] _04110_ _04874_ _04876_ vssd1 vssd1 vccd1
+ vccd1 _04878_ sky130_fd_sc_hd__mux4_1
XFILLER_108_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11123_ rbzero.texV\[5\] _03841_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__xor2_1
XFILLER_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16980_ _09398_ _09401_ _09519_ vssd1 vssd1 vccd1 vccd1 _09521_ sky130_fd_sc_hd__and3_1
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15931_ _07623_ _07920_ _07919_ vssd1 vssd1 vccd1 vccd1 _08545_ sky130_fd_sc_hd__o21bai_1
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11054_ _03780_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__buf_2
XFILLER_89_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18650_ rbzero.debug_overlay.vplaneY\[-6\] rbzero.wall_tracer.rayAddendY\[-6\] _02381_
+ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__o21ai_1
XFILLER_231_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15862_ _07689_ _07819_ _07690_ _08475_ vssd1 vssd1 vccd1 vccd1 _08476_ sky130_fd_sc_hd__a31o_1
XFILLER_190_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17601_ _10136_ _10137_ vssd1 vssd1 vccd1 vccd1 _10138_ sky130_fd_sc_hd__nor2_1
XFILLER_225_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14813_ rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__xor2_1
XFILLER_218_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18581_ _02320_ _02321_ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__xnor2_1
X_15793_ _08380_ _08375_ _08379_ vssd1 vssd1 vccd1 vccd1 _08407_ sky130_fd_sc_hd__and3_1
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17532_ _10055_ _10067_ vssd1 vssd1 vccd1 vccd1 _10069_ sky130_fd_sc_hd__or2_1
XFILLER_40_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14744_ rbzero.debug_overlay.playerY\[-6\] _07357_ vssd1 vssd1 vccd1 vccd1 _07358_
+ sky130_fd_sc_hd__or2_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ net17 net18 vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__nor2_1
XFILLER_233_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_146 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_146/HI o_rgb[4] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_157 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_157/HI o_rgb[19]
+ sky130_fd_sc_hd__conb_1
XFILLER_225_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17463_ _09999_ _10000_ vssd1 vssd1 vccd1 vccd1 _10001_ sky130_fd_sc_hd__or2_1
XFILLER_205_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10907_ rbzero.tex_b0\[44\] rbzero.tex_b0\[43\] _03671_ vssd1 vssd1 vccd1 vccd1 _03680_
+ sky130_fd_sc_hd__mux2_1
XFILLER_232_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14675_ _07311_ vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11887_ rbzero.row_render.texu\[5\] rbzero.row_render.texu\[4\] rbzero.row_render.texu\[3\]
+ rbzero.row_render.texu\[2\] _03288_ _04592_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__mux4_1
XFILLER_233_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19202_ rbzero.spi_registers.new_vshift\[4\] _02775_ vssd1 vssd1 vccd1 vccd1 _02781_
+ sky130_fd_sc_hd__or2_1
X_16414_ _09021_ _09023_ vssd1 vssd1 vccd1 vccd1 _09024_ sky130_fd_sc_hd__and2_1
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13626_ _06310_ _06312_ _06314_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__o21a_1
X_10838_ rbzero.tex_g0\[13\] rbzero.tex_g0\[12\] _03638_ vssd1 vssd1 vccd1 vccd1 _03644_
+ sky130_fd_sc_hd__mux2_1
X_17394_ _09930_ _09931_ vssd1 vssd1 vccd1 vccd1 _09932_ sky130_fd_sc_hd__and2_1
XFILLER_220_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19133_ rbzero.othery\[3\] _02723_ _02736_ _02728_ vssd1 vssd1 vccd1 vccd1 _00740_
+ sky130_fd_sc_hd__o211a_1
X_16345_ _08953_ _08954_ vssd1 vssd1 vccd1 vccd1 _08956_ sky130_fd_sc_hd__nand2_1
XFILLER_160_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13557_ _06204_ _06245_ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__xor2_1
X_10769_ rbzero.tex_g0\[46\] rbzero.tex_g0\[45\] _03605_ vssd1 vssd1 vccd1 vccd1 _03608_
+ sky130_fd_sc_hd__mux2_1
XFILLER_121_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12508_ rbzero.wall_tracer.visualWallDist\[3\] _05190_ _03789_ vssd1 vssd1 vccd1
+ vccd1 _05197_ sky130_fd_sc_hd__a21o_1
X_19064_ _02694_ vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__clkbuf_1
X_16276_ _07742_ _07591_ _07520_ _08135_ vssd1 vssd1 vccd1 vccd1 _08887_ sky130_fd_sc_hd__a2bb2o_1
X_13488_ _05839_ _05878_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__nand2_1
XFILLER_199_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18015_ _01758_ _01796_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15227_ _04935_ _07664_ vssd1 vssd1 vccd1 vccd1 _07841_ sky130_fd_sc_hd__or2_1
X_12439_ _05130_ vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15158_ _07764_ _07770_ _07771_ vssd1 vssd1 vccd1 vccd1 _07772_ sky130_fd_sc_hd__a21oi_1
XFILLER_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14109_ _05641_ _06321_ vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__and2_1
X_15089_ _07195_ _07198_ _07213_ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__o21a_1
X_19966_ _03119_ vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__clkinv_2
Xfanout109 net115 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__buf_2
XFILLER_141_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18917_ rbzero.pov.spi_buffer\[8\] rbzero.pov.ready_buffer\[8\] _02608_ vssd1 vssd1
+ vccd1 vccd1 _02617_ sky130_fd_sc_hd__mux2_1
XFILLER_171_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19897_ _03112_ vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__clkinv_2
XFILLER_41_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18848_ _02563_ _02564_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__nand2_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18779_ _02428_ rbzero.debug_overlay.vplaneY\[-4\] _02498_ _02499_ vssd1 vssd1 vccd1
+ vccd1 _02501_ sky130_fd_sc_hd__nor4_1
XFILLER_209_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20810_ _00028_ _00826_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20741_ net107 _00757_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20672_ net70 _00688_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21224_ _00273_ _01240_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21155_ _00204_ _01171_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20106_ _09245_ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__buf_2
XFILLER_137_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21086_ _00135_ _01102_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20037_ _03125_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__clkbuf_8
XFILLER_86_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ rbzero.tex_b1\[53\] rbzero.tex_b1\[52\] _04032_ vssd1 vssd1 vccd1 vccd1 _04524_
+ sky130_fd_sc_hd__mux2_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _05475_ _05476_ _05478_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__mux2_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11741_ rbzero.tex_b0\[49\] rbzero.tex_b0\[48\] _04013_ vssd1 vssd1 vccd1 vccd1 _04456_
+ sky130_fd_sc_hd__mux2_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20939_ net100 _00955_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ss_buffer\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14460_ _07102_ _07146_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__nand2_1
XFILLER_159_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ rbzero.tex_g1\[22\] _04374_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__and2_1
XFILLER_241_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13411_ _06073_ _06074_ _06080_ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__a21o_1
X_10623_ _03531_ vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__clkbuf_1
X_14391_ _07007_ _07078_ _07079_ _07049_ vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_224_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16130_ _08739_ _08740_ vssd1 vssd1 vccd1 vccd1 _08742_ sky130_fd_sc_hd__and2_1
XFILLER_195_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13342_ _05626_ _06010_ _05715_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10554_ rbzero.tex_r0\[20\] rbzero.tex_r0\[19\] _03490_ vssd1 vssd1 vccd1 vccd1 _03495_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16061_ _07788_ _07916_ vssd1 vssd1 vccd1 vccd1 _08674_ sky130_fd_sc_hd__nor2_1
X_13273_ _05956_ _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__xor2_1
XFILLER_108_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10485_ rbzero.tex_r0\[53\] rbzero.tex_r0\[52\] _03457_ vssd1 vssd1 vccd1 vccd1 _03459_
+ sky130_fd_sc_hd__mux2_1
XFILLER_237_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15012_ _07616_ _07619_ _07618_ _07625_ vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__o22a_1
X_12224_ o_vsync rbzero.wall_tracer.state\[9\] _03292_ vssd1 vssd1 vccd1 vccd1 _04924_
+ sky130_fd_sc_hd__and3_1
XFILLER_154_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19820_ _03105_ vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__clkinv_2
XFILLER_68_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ net52 _04825_ net27 vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__and3_1
XFILLER_64_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11106_ _03820_ _03822_ _03824_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__or3b_2
XFILLER_111_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19751_ rbzero.pov.ready_buffer\[1\] _03069_ _03070_ rbzero.debug_overlay.vplaneY\[-8\]
+ _02832_ vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__o221a_1
X_16963_ _09501_ _09503_ vssd1 vssd1 vccd1 vccd1 _09505_ sky130_fd_sc_hd__and2_1
X_12086_ net26 _04793_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__nand2_1
XFILLER_238_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18702_ _02428_ rbzero.wall_tracer.rayAddendY\[0\] vssd1 vssd1 vccd1 vccd1 _02429_
+ sky130_fd_sc_hd__nor2_1
XFILLER_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15914_ _07873_ _07904_ vssd1 vssd1 vccd1 vccd1 _08528_ sky130_fd_sc_hd__and2_1
X_11037_ rbzero.otherx\[0\] _03742_ _03746_ rbzero.otherx\[3\] vssd1 vssd1 vccd1 vccd1
+ _03765_ sky130_fd_sc_hd__a22o_1
XFILLER_209_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19682_ rbzero.debug_overlay.playerY\[1\] _03032_ rbzero.debug_overlay.playerY\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__o21ai_1
X_16894_ _09172_ _09434_ _09435_ _09170_ vssd1 vssd1 vccd1 vccd1 _09436_ sky130_fd_sc_hd__a22o_1
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18633_ _03746_ _07491_ _02365_ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__a21oi_1
XFILLER_225_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15845_ _08110_ _08171_ _08457_ _08458_ vssd1 vssd1 vccd1 vccd1 _08459_ sky130_fd_sc_hd__a31o_2
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18564_ _02274_ _02191_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__and2_1
XFILLER_206_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15776_ _08368_ _08389_ vssd1 vssd1 vccd1 vccd1 _08390_ sky130_fd_sc_hd__xnor2_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12988_ _05670_ _05676_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__and2b_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17515_ _09022_ _08890_ _08851_ _08979_ vssd1 vssd1 vccd1 vccd1 _10052_ sky130_fd_sc_hd__or4_1
XFILLER_205_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14727_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__buf_2
XFILLER_75_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18495_ _02226_ _02240_ _02236_ _03818_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__a31o_1
X_11939_ _04630_ net11 _04646_ _04649_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__a31o_1
XFILLER_233_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17446_ _09981_ _09982_ _09977_ vssd1 vssd1 vccd1 vccd1 _09984_ sky130_fd_sc_hd__a21o_1
XFILLER_33_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14658_ rbzero.wall_tracer.trackDistX\[9\] rbzero.wall_tracer.trackDistY\[9\] _05025_
+ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__mux2_1
XFILLER_162_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13609_ _06277_ _06296_ _06297_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__a21bo_1
XFILLER_92_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17377_ _08890_ _08850_ _08979_ _08596_ vssd1 vssd1 vccd1 vccd1 _09915_ sky130_fd_sc_hd__o22a_1
XFILLER_158_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14589_ _07252_ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__clkbuf_4
XFILLER_159_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19116_ _02727_ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__clkbuf_4
X_16328_ _08792_ _08801_ _08938_ vssd1 vssd1 vccd1 vccd1 _08939_ sky130_fd_sc_hd__a21o_1
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19047_ rbzero.pov.spi_buffer\[70\] rbzero.pov.ready_buffer\[70\] _02607_ vssd1 vssd1
+ vccd1 vccd1 _02685_ sky130_fd_sc_hd__mux2_1
XFILLER_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16259_ _08864_ _08869_ vssd1 vssd1 vccd1 vccd1 _08870_ sky130_fd_sc_hd__xnor2_1
XFILLER_199_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19949_ _03118_ vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__clkinv_2
XFILLER_228_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20724_ net94 _00740_ vssd1 vssd1 vccd1 vccd1 rbzero.othery\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20655_ net63 _00671_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20586_ net95 _00602_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10270_ _03343_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21207_ _00256_ _01223_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21138_ _00187_ _01154_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13960_ _06310_ _06423_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__nor2_1
XFILLER_150_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21069_ _00118_ _01085_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12911_ _05505_ _05430_ _05599_ _05586_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__a211o_1
XFILLER_207_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13891_ _06578_ _06579_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__xnor2_1
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15630_ _08231_ _08239_ _08243_ vssd1 vssd1 vccd1 vccd1 _08244_ sky130_fd_sc_hd__o21a_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12842_ _05399_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__buf_2
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _08086_ _07970_ _07554_ _07697_ vssd1 vssd1 vccd1 vccd1 _08175_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _05452_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__clkbuf_4
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17300_ _08760_ _08780_ vssd1 vssd1 vccd1 vccd1 _09839_ sky130_fd_sc_hd__nor2_1
XFILLER_163_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14512_ _07102_ _07191_ vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__nand2_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18280_ _09279_ _02050_ _02001_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__a21o_1
XFILLER_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _04323_ _04437_ _04438_ _04439_ _03972_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__o221a_1
XFILLER_202_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15492_ _08074_ _08105_ vssd1 vssd1 vccd1 vccd1 _08106_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _09766_ _09767_ _09768_ vssd1 vssd1 vccd1 vccd1 _09771_ sky130_fd_sc_hd__a21o_1
X_14443_ _07039_ _07047_ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__or2_1
XFILLER_70_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11655_ _04370_ _04371_ _04099_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__mux2_1
XFILLER_230_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout80 net83 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__buf_2
XFILLER_243_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout91 net92 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17162_ _09163_ _07837_ _09700_ vssd1 vssd1 vccd1 vccd1 _09702_ sky130_fd_sc_hd__a21o_1
XFILLER_7_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10606_ _03522_ vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14374_ _05408_ _07057_ _07062_ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__a21oi_1
XFILLER_161_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11586_ rbzero.tex_g0\[19\] rbzero.tex_g0\[18\] _04119_ vssd1 vssd1 vccd1 vccd1 _04303_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16113_ _08724_ vssd1 vssd1 vccd1 vccd1 _08725_ sky130_fd_sc_hd__clkbuf_4
XFILLER_196_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13325_ _05999_ _06013_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__xor2_1
XFILLER_128_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10537_ rbzero.tex_r0\[28\] rbzero.tex_r0\[27\] _03479_ vssd1 vssd1 vccd1 vccd1 _03486_
+ sky130_fd_sc_hd__mux2_1
X_17093_ _09631_ _09633_ vssd1 vssd1 vccd1 vccd1 _09634_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16044_ _08502_ _08524_ _08501_ vssd1 vssd1 vccd1 vccd1 _08657_ sky130_fd_sc_hd__a21boi_1
XFILLER_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13256_ _05896_ _05941_ _05942_ _05944_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__a22o_1
X_10468_ rbzero.tex_r0\[61\] rbzero.tex_r0\[60\] _03446_ vssd1 vssd1 vccd1 vccd1 _03450_
+ sky130_fd_sc_hd__mux2_1
XFILLER_100_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _04873_ _04874_ gpout5.clk_div\[0\] _04912_ vssd1 vssd1 vccd1 vccd1 _04913_
+ sky130_fd_sc_hd__a31o_1
X_13187_ _05765_ _05777_ _05875_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__a21oi_1
XFILLER_83_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10399_ rbzero.tex_r1\[27\] rbzero.tex_r1\[28\] _03411_ vssd1 vssd1 vccd1 vccd1 _03412_
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12138_ net30 net31 _04844_ net32 vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__a22oi_1
X_19803_ _04113_ _03096_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__nand2_1
XFILLER_170_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17995_ _01766_ _01776_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__nand2_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16946_ _09485_ _09487_ vssd1 vssd1 vccd1 vccd1 _09488_ sky130_fd_sc_hd__xnor2_1
X_12069_ _04768_ o_rgb[23] _04775_ _04776_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__a211o_1
XFILLER_111_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19734_ _03062_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__buf_2
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19665_ rbzero.pov.ready_buffer\[51\] _02836_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__nand2_1
XFILLER_237_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16877_ _09403_ _09418_ vssd1 vssd1 vccd1 vccd1 _09419_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18616_ rbzero.map_rom.f3 _02351_ _09274_ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__mux2_1
X_15828_ _08413_ _08439_ vssd1 vssd1 vccd1 vccd1 _08442_ sky130_fd_sc_hd__nand2_1
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19596_ rbzero.pov.ready_buffer\[65\] _07539_ _02962_ vssd1 vssd1 vccd1 vccd1 _02974_
+ sky130_fd_sc_hd__mux2_1
XFILLER_231_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18547_ _02277_ _02280_ _02288_ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a21o_1
XFILLER_234_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15759_ _08365_ _08367_ _08371_ vssd1 vssd1 vccd1 vccd1 _08373_ sky130_fd_sc_hd__nor3_1
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18478_ _02212_ _02215_ _02225_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a21o_1
XFILLER_166_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17429_ _09965_ _09966_ vssd1 vssd1 vccd1 vccd1 _09967_ sky130_fd_sc_hd__xor2_1
XFILLER_127_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20440_ net138 _00471_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20371_ net92 _00404_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.a6 sky130_fd_sc_hd__dfxtp_2
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20707_ net99 _00723_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11440_ rbzero.tex_r1\[19\] rbzero.tex_r1\[18\] _04000_ vssd1 vssd1 vccd1 vccd1 _04158_
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20638_ net55 _00654_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11371_ gpout0.hpos\[3\] _04082_ _04084_ gpout0.hpos\[2\] _04089_ vssd1 vssd1 vccd1
+ vccd1 _04090_ sky130_fd_sc_hd__o221a_1
X_20569_ net139 _00585_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_164_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13110_ _05792_ _05794_ _05798_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__or3_1
X_10322_ rbzero.tex_r1\[63\] net48 _03366_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__mux2_1
X_14090_ _06752_ _06778_ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__xnor2_1
XFILLER_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13041_ _05715_ _05728_ _05726_ _05607_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__o22ai_1
XFILLER_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10253_ rbzero.tex_b1\[32\] rbzero.tex_b1\[33\] _03333_ vssd1 vssd1 vccd1 vccd1 _03335_
+ sky130_fd_sc_hd__mux2_1
XFILLER_106_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10184_ _03294_ _03296_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__nor2_1
XFILLER_26_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16800_ _04940_ vssd1 vssd1 vccd1 vccd1 _09345_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17780_ _01525_ _01563_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__xnor2_2
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14992_ _07507_ _07542_ _07549_ _07575_ vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__or4_1
XFILLER_8_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16731_ rbzero.wall_tracer.trackDistX\[-12\] _09276_ _09278_ _09284_ vssd1 vssd1
+ vccd1 vccd1 _00541_ sky130_fd_sc_hd__o22a_1
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13943_ _06625_ _06623_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__xor2_1
XFILLER_208_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19450_ rbzero.pov.spi_buffer\[22\] rbzero.pov.spi_buffer\[23\] _02888_ vssd1 vssd1
+ vccd1 vccd1 _02892_ sky130_fd_sc_hd__mux2_1
XFILLER_207_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16662_ _09257_ vssd1 vssd1 vccd1 vccd1 _09259_ sky130_fd_sc_hd__buf_2
XFILLER_234_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13874_ _06504_ _06562_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__nand2_1
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18401_ rbzero.debug_overlay.vplaneX\[-6\] rbzero.wall_tracer.rayAddendX\[-6\] _02154_
+ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__o21ai_1
X_15613_ _07467_ _07508_ vssd1 vssd1 vccd1 vccd1 _08227_ sky130_fd_sc_hd__nor2_1
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12825_ _05513_ _05472_ _05462_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__mux2_2
X_19381_ _02860_ vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__clkinv_2
X_16593_ _09052_ _09201_ vssd1 vssd1 vccd1 vccd1 _09202_ sky130_fd_sc_hd__and2_1
XFILLER_216_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18332_ rbzero.wall_tracer.trackDistY\[4\] rbzero.wall_tracer.stepDistY\[4\] vssd1
+ vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__nor2_1
X_15544_ _08152_ _08157_ vssd1 vssd1 vccd1 vccd1 _08158_ sky130_fd_sc_hd__xnor2_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12756_ _05444_ _05428_ _05399_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__a21o_1
XFILLER_128_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18263_ _02033_ _02034_ _02035_ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__or3_1
XFILLER_124_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11707_ rbzero.tex_g1\[53\] rbzero.tex_g1\[52\] _04378_ vssd1 vssd1 vccd1 vccd1 _04423_
+ sky130_fd_sc_hd__mux2_1
XFILLER_188_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15475_ _08084_ _08087_ _08088_ vssd1 vssd1 vccd1 vccd1 _08089_ sky130_fd_sc_hd__a21o_1
XFILLER_128_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12687_ _05373_ _05375_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__or2_1
X_17214_ _09526_ _09630_ _09753_ vssd1 vssd1 vccd1 vccd1 _09754_ sky130_fd_sc_hd__a21oi_1
XFILLER_129_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14426_ _05517_ _05499_ vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__nor2_1
XFILLER_129_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18194_ _01932_ _01973_ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__xnor2_1
XFILLER_198_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11638_ _04353_ _04354_ _04014_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__mux2_1
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17145_ _09684_ _08735_ vssd1 vssd1 vccd1 vccd1 _09685_ sky130_fd_sc_hd__nor2_1
X_14357_ _05431_ _07024_ vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__nor2_1
XFILLER_144_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11569_ _04280_ _04281_ _04283_ _04286_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__or4_1
XFILLER_156_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13308_ _05984_ _05988_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__xor2_1
XFILLER_143_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17076_ _09469_ _09480_ _09616_ vssd1 vssd1 vccd1 vccd1 _09617_ sky130_fd_sc_hd__a21bo_1
XFILLER_196_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14288_ _06453_ _06402_ _06976_ vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__o21ai_1
XFILLER_170_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16027_ _07519_ rbzero.wall_tracer.stepDistX\[4\] vssd1 vssd1 vccd1 vccd1 _08640_
+ sky130_fd_sc_hd__nand2_2
XFILLER_143_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13239_ _05906_ _05924_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__nor2_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17978_ _01629_ _01643_ _01759_ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__a21bo_1
XFILLER_211_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16929_ _08923_ _09470_ _07835_ vssd1 vssd1 vccd1 vccd1 _09471_ sky130_fd_sc_hd__a21o_1
X_19717_ rbzero.pov.ready_buffer\[38\] _03056_ _03059_ rbzero.debug_overlay.facingX\[-4\]
+ _03065_ vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__o221a_1
XFILLER_211_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19648_ _08574_ _03008_ _03014_ _03015_ vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__a211oi_1
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19579_ _02740_ _02833_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__nor2_4
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20423_ net126 _00454_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20354_ gpout2.clk_div\[0\] gpout2.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__nand2_1
XFILLER_122_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20285_ _03257_ vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__clkinv_2
XTAP_6206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10940_ _03697_ vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10871_ _03661_ vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12610_ _05277_ _05289_ _05296_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__o21a_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13590_ _06277_ _06278_ vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__nor2_1
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ _05155_ _05158_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__xnor2_2
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15260_ _07869_ _07870_ _07872_ vssd1 vssd1 vccd1 vccd1 _07874_ sky130_fd_sc_hd__a21o_1
XFILLER_200_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12472_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] vssd1
+ vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__and2_1
XFILLER_32_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14211_ _06887_ _06897_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__xnor2_1
XFILLER_240_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11423_ rbzero.tex_r1\[40\] _03959_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__and2_1
X_15191_ _07567_ vssd1 vssd1 vccd1 vccd1 _07805_ sky130_fd_sc_hd__clkbuf_4
XFILLER_126_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14142_ _06829_ _06830_ vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__and2_1
X_11354_ _03290_ _04072_ _04071_ _03293_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__a22o_1
XFILLER_180_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10305_ rbzero.tex_b1\[7\] rbzero.tex_b1\[8\] _03355_ vssd1 vssd1 vccd1 vccd1 _03362_
+ sky130_fd_sc_hd__mux2_1
XFILLER_180_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14073_ _05668_ _06321_ vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__nand2_1
XFILLER_152_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11285_ _03932_ _03999_ _04002_ _04003_ _03923_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__o221a_1
X_18950_ _02634_ vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__clkbuf_1
X_17901_ _01649_ _01683_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__xnor2_1
X_13024_ _05612_ _05700_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__nand2_1
X_10236_ rbzero.tex_b1\[40\] rbzero.tex_b1\[41\] _03322_ vssd1 vssd1 vccd1 vccd1 _03326_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18881_ rbzero.spi_registers.spi_counter\[2\] rbzero.spi_registers.spi_counter\[1\]
+ rbzero.spi_registers.spi_counter\[0\] _02576_ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__and4_1
XTAP_6740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17832_ _01613_ _01614_ _01615_ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__a21oi_1
XTAP_6773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17763_ _01545_ _01546_ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__and2_1
X_14975_ _07476_ _07490_ _07587_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__nand3_1
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19502_ rbzero.pov.spi_buffer\[47\] rbzero.pov.spi_buffer\[48\] _02910_ vssd1 vssd1
+ vccd1 vccd1 _02919_ sky130_fd_sc_hd__mux2_1
X_16714_ rbzero.wall_tracer.wall\[0\] rbzero.row_render.wall\[0\] _09269_ vssd1 vssd1
+ vccd1 vccd1 _09270_ sky130_fd_sc_hd__mux2_1
XFILLER_212_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13926_ _06610_ _06613_ vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__and2b_1
X_17694_ _01476_ _01477_ _01471_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__a21o_1
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19433_ rbzero.pov.spi_buffer\[14\] rbzero.pov.spi_buffer\[15\] _02877_ vssd1 vssd1
+ vccd1 vccd1 _02883_ sky130_fd_sc_hd__mux2_1
X_16645_ _04198_ _09244_ vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__nor2_1
XFILLER_62_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13857_ _06479_ _06539_ _06545_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__o21a_1
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12808_ _05453_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__buf_2
X_19364_ _02859_ vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__clkinv_2
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16576_ _08398_ _09051_ _09048_ vssd1 vssd1 vccd1 vccd1 _09185_ sky130_fd_sc_hd__o21a_1
X_13788_ _06467_ _06475_ _06476_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__a21boi_1
XFILLER_222_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18315_ _01997_ _02079_ _02080_ _02013_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__a31o_1
XFILLER_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15527_ _08135_ _08136_ _08139_ _08140_ vssd1 vssd1 vccd1 vccd1 _08141_ sky130_fd_sc_hd__a31oi_2
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12739_ _05427_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__clkbuf_2
XFILLER_31_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19295_ _04920_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__clkbuf_4
XFILLER_148_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18246_ rbzero.wall_tracer.trackDistY\[-8\] rbzero.wall_tracer.stepDistY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__nor2_1
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15458_ _08053_ _08055_ _08071_ vssd1 vssd1 vccd1 vccd1 _08072_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14409_ _07080_ _07083_ _07090_ _07097_ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__o31ai_4
X_18177_ _10095_ _08985_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__nor2_1
XFILLER_239_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ _07955_ _07957_ vssd1 vssd1 vccd1 vccd1 _08003_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17128_ _09022_ _08718_ _08855_ _08750_ vssd1 vssd1 vccd1 vccd1 _09668_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_237_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17059_ _09598_ _09599_ vssd1 vssd1 vccd1 vccd1 _09600_ sky130_fd_sc_hd__nor2_1
XFILLER_239_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20070_ _03125_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__buf_6
XFILLER_83_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20972_ net70 _00988_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20406_ net128 _00437_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_107_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21386_ net109 _01402_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20337_ _02146_ _02152_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__and2b_1
XFILLER_134_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11070_ _03793_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__clkbuf_4
XFILLER_153_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20268_ _03255_ vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__clkinv_2
XTAP_6036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20199_ rbzero.texV\[4\] _03137_ _03142_ _03220_ vssd1 vssd1 vccd1 vccd1 _01322_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _05196_ _07368_ _07373_ _05186_ vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__a31oi_4
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ net17 _04677_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__nor2_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13711_ _06372_ _06399_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__or2_1
XFILLER_245_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10923_ _03688_ vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14691_ rbzero.wall_tracer.stepDistX\[0\] _07202_ _07316_ vssd1 vssd1 vccd1 vccd1
+ _07320_ sky130_fd_sc_hd__mux2_1
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16430_ _08771_ _08788_ _09037_ _09038_ _09039_ vssd1 vssd1 vccd1 vccd1 _09040_ sky130_fd_sc_hd__a32o_1
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13642_ _06330_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__buf_2
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10854_ _03652_ vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _08859_ _08860_ _08970_ vssd1 vssd1 vccd1 vccd1 _08971_ sky130_fd_sc_hd__o21a_1
XFILLER_201_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13573_ _06214_ _06254_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__nand2_2
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _03604_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__clkbuf_4
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18100_ _01879_ _01880_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__and2_1
XFILLER_125_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _07924_ _07925_ vssd1 vssd1 vccd1 vccd1 _07926_ sky130_fd_sc_hd__nor2_1
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12524_ _03815_ _05076_ _05077_ _05212_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__a31o_1
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19080_ rbzero.spi_registers.spi_counter\[3\] rbzero.spi_registers.spi_counter\[2\]
+ _02577_ _02702_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__or4_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _08883_ _08902_ vssd1 vssd1 vccd1 vccd1 _08903_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18031_ _01690_ _01701_ _01688_ vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15243_ _07852_ _07853_ _07855_ vssd1 vssd1 vccd1 vccd1 _07857_ sky130_fd_sc_hd__a21o_1
XFILLER_201_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12455_ rbzero.debug_overlay.facingX\[0\] rbzero.wall_tracer.rayAddendX\[8\] vssd1
+ vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__or2_1
XFILLER_138_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11406_ rbzero.tex_r1\[53\] rbzero.tex_r1\[52\] _04119_ vssd1 vssd1 vccd1 vccd1 _04124_
+ sky130_fd_sc_hd__mux2_1
X_15174_ _07517_ vssd1 vssd1 vccd1 vccd1 _07788_ sky130_fd_sc_hd__clkbuf_4
X_12386_ _05056_ _05058_ _05064_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__a21oi_1
XFILLER_181_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14125_ _06761_ _06770_ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__xnor2_1
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11337_ rbzero.row_render.size\[1\] vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__inv_2
XFILLER_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19982_ _03121_ vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__clkinv_2
XFILLER_158_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14056_ _06700_ _06743_ _06744_ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__a21oi_1
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18933_ _02625_ vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11268_ rbzero.tex_r0\[19\] rbzero.tex_r0\[18\] _03974_ vssd1 vssd1 vccd1 vccd1 _03987_
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ _05667_ _05686_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__and2_1
XFILLER_122_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10219_ rbzero.tex_b1\[48\] rbzero.tex_b1\[49\] _03311_ vssd1 vssd1 vccd1 vccd1 _03317_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18864_ rbzero.spi_registers.spi_cmd\[2\] _02578_ rbzero.spi_registers.spi_cmd\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__a21o_1
X_11199_ _03863_ _03852_ _03860_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__nor3_1
XTAP_6570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17815_ _01564_ _01598_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18795_ _02516_ vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__clkbuf_1
XTAP_5880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17746_ _09166_ _08851_ _08979_ _09684_ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__o22a_1
XFILLER_36_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14958_ _07408_ rbzero.wall_tracer.stepDistY\[-8\] _07352_ vssd1 vssd1 vccd1 vccd1
+ _07572_ sky130_fd_sc_hd__a21oi_4
XFILLER_78_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13909_ _06528_ _06594_ _06595_ _06597_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__a22oi_2
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17677_ _01459_ _01461_ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__and2b_1
XFILLER_63_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14889_ _07341_ _05096_ _07336_ vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__o21a_1
XFILLER_36_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16628_ _09234_ _09236_ vssd1 vssd1 vccd1 vccd1 _09237_ sky130_fd_sc_hd__xor2_4
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19416_ rbzero.pov.spi_buffer\[6\] rbzero.pov.spi_buffer\[7\] _02866_ vssd1 vssd1
+ vccd1 vccd1 _02874_ sky130_fd_sc_hd__mux2_1
XFILLER_211_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16559_ _09165_ _09167_ vssd1 vssd1 vccd1 vccd1 _09168_ sky130_fd_sc_hd__xnor2_1
X_19347_ _02857_ vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__clkinv_2
XFILLER_204_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19278_ _02823_ vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18229_ _01997_ _02005_ _02006_ _02001_ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__a31o_1
XFILLER_163_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21240_ _00289_ _01256_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21171_ _00220_ _01187_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20122_ _03153_ _03154_ _03155_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__o21ai_1
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20053_ _03128_ vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__clkinv_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20955_ net91 _00971_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ net66 _00902_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10570_ _03503_ vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12240_ rbzero.debug_overlay.playerY\[0\] _03743_ _03798_ vssd1 vssd1 vccd1 vccd1
+ _04934_ sky130_fd_sc_hd__mux2_1
XFILLER_147_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12171_ _04591_ _04080_ _04628_ _04101_ _04874_ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_
+ sky130_fd_sc_hd__mux4_1
XFILLER_68_1346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21369_ _00392_ _01385_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11122_ _03838_ _03837_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__nand2_1
XFILLER_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15930_ _08534_ _08543_ vssd1 vssd1 vccd1 vccd1 _08544_ sky130_fd_sc_hd__xnor2_1
X_11053_ gpout0.hpos\[5\] vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__buf_2
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15861_ _07223_ _07096_ _07101_ _07224_ vssd1 vssd1 vccd1 vccd1 _08475_ sky130_fd_sc_hd__o211a_1
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17600_ _10133_ _10135_ vssd1 vssd1 vccd1 vccd1 _10137_ sky130_fd_sc_hd__and2_1
XTAP_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ _07403_ _07425_ vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__xnor2_1
XTAP_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18580_ _02299_ _02304_ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__nand2_1
X_15792_ _08399_ _08405_ vssd1 vssd1 vccd1 vccd1 _08406_ sky130_fd_sc_hd__nor2_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _10055_ _10067_ vssd1 vssd1 vccd1 vccd1 _10068_ sky130_fd_sc_hd__nand2_1
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14743_ rbzero.debug_overlay.playerY\[-7\] rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerY\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__or3_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ net15 vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__buf_2
XFILLER_45_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17462_ _09997_ _09998_ _09973_ vssd1 vssd1 vccd1 vccd1 _10000_ sky130_fd_sc_hd__a21oi_1
XFILLER_233_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_147 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_147/HI o_rgb[5] sky130_fd_sc_hd__conb_1
X_10906_ _03679_ vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__clkbuf_1
Xtop_ew_algofoogle_158 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_158/HI o_rgb[20]
+ sky130_fd_sc_hd__conb_1
XFILLER_229_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14674_ rbzero.wall_tracer.stepDistX\[-8\] _07165_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _07311_ sky130_fd_sc_hd__mux2_1
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11886_ _04591_ _04598_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__or2_1
X_16413_ _09022_ _07886_ _09020_ vssd1 vssd1 vccd1 vccd1 _09023_ sky130_fd_sc_hd__o21ai_1
X_19201_ rbzero.spi_registers.vshift\[3\] _02774_ _02779_ _02780_ vssd1 vssd1 vccd1
+ vccd1 _00764_ sky130_fd_sc_hd__o211a_1
X_13625_ _06313_ _06305_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__or2b_1
XFILLER_232_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17393_ _09919_ _09929_ vssd1 vssd1 vccd1 vccd1 _09931_ sky130_fd_sc_hd__or2_1
XFILLER_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10837_ _03643_ vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19132_ rbzero.spi_registers.new_other\[3\] _02725_ vssd1 vssd1 vccd1 vccd1 _02736_
+ sky130_fd_sc_hd__or2_1
X_16344_ _08953_ _08954_ vssd1 vssd1 vccd1 vccd1 _08955_ sky130_fd_sc_hd__or2_2
XFILLER_164_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13556_ _06237_ _06244_ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__xor2_1
XFILLER_160_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10768_ _03607_ vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12507_ _05184_ _05195_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__xor2_2
XFILLER_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19063_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.spi_buffer\[2\]
+ _02690_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__mux2_1
X_16275_ _07742_ _08223_ _07591_ _07790_ vssd1 vssd1 vccd1 vccd1 _08886_ sky130_fd_sc_hd__or4_1
XFILLER_199_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13487_ _06165_ _06175_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__or2_2
XFILLER_173_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10699_ rbzero.tex_g1\[14\] rbzero.tex_g1\[15\] _03563_ vssd1 vssd1 vccd1 vccd1 _03571_
+ sky130_fd_sc_hd__mux2_1
XFILLER_218_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18014_ _01760_ _01795_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__xnor2_1
XFILLER_199_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15226_ _07686_ _07695_ vssd1 vssd1 vccd1 vccd1 _07840_ sky130_fd_sc_hd__nor2_2
XFILLER_145_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12438_ _05129_ _03733_ _05028_ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__mux2_1
XFILLER_126_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15157_ _07758_ _07763_ vssd1 vssd1 vccd1 vccd1 _07771_ sky130_fd_sc_hd__nor2_1
XFILLER_154_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12369_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[9\] vssd1
+ vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__or2_1
XFILLER_181_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14108_ _06777_ _06776_ _06754_ vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__a21o_1
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15088_ rbzero.wall_tracer.stepDistY\[-1\] vssd1 vssd1 vccd1 vccd1 _07702_ sky130_fd_sc_hd__inv_2
X_19965_ _03119_ vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__clkinv_2
XFILLER_102_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14039_ _06712_ _06726_ _06727_ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__a21bo_1
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18916_ _02616_ vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__clkbuf_1
XTAP_7090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19896_ _03112_ vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__clkinv_2
XFILLER_110_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18847_ _02510_ rbzero.wall_tracer.rayAddendY\[10\] vssd1 vssd1 vccd1 vccd1 _02564_
+ sky130_fd_sc_hd__xor2_1
XFILLER_68_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18778_ _02428_ rbzero.debug_overlay.vplaneY\[-4\] _02498_ _02499_ vssd1 vssd1 vccd1
+ vccd1 _02500_ sky130_fd_sc_hd__o22a_1
XFILLER_227_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17729_ _01494_ _01495_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__or2_1
XFILLER_247_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20740_ net105 _00756_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20671_ net74 _00687_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21223_ _00272_ _01239_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21154_ _00203_ _01170_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20105_ _03093_ _03140_ _03141_ _03137_ rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1
+ _01307_ sky130_fd_sc_hd__a32o_1
XFILLER_28_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21085_ _00134_ _01101_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20036_ _03126_ vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__clkinv_2
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _04007_ _04450_ _04454_ _03956_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__a211o_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ net87 _00954_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.mosi sky130_fd_sc_hd__dfxtp_1
XFILLER_230_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ rbzero.tex_g1\[21\] rbzero.tex_g1\[20\] _04378_ vssd1 vssd1 vccd1 vccd1 _04387_
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20869_ net54 _00885_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13410_ _06073_ _06074_ _06080_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__nand3_1
XFILLER_35_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10622_ rbzero.tex_g1\[51\] rbzero.tex_g1\[52\] _03530_ vssd1 vssd1 vccd1 vccd1 _03531_
+ sky130_fd_sc_hd__mux2_1
X_14390_ _07029_ _05404_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__and2_1
XFILLER_122_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13341_ _05986_ _05987_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__xor2_1
XFILLER_127_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10553_ _03494_ vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16060_ _08669_ _08672_ vssd1 vssd1 vccd1 vccd1 _08673_ sky130_fd_sc_hd__nand2_1
XFILLER_127_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13272_ _05914_ _05957_ _05958_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__o22a_1
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10484_ _03458_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15011_ _07624_ vssd1 vssd1 vccd1 vccd1 _07625_ sky130_fd_sc_hd__buf_2
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12223_ _03791_ _03730_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__nor2_1
XFILLER_123_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12154_ _04115_ _04859_ _04860_ gpout4.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _04861_
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11105_ gpout0.hpos\[7\] gpout0.hpos\[8\] _03823_ gpout0.hpos\[9\] vssd1 vssd1 vccd1
+ vccd1 _03824_ sky130_fd_sc_hd__a31o_1
XFILLER_46_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19750_ rbzero.pov.ready_buffer\[0\] _03067_ _03068_ rbzero.debug_overlay.vplaneY\[-9\]
+ _03015_ vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__a221o_1
XFILLER_231_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16962_ _09501_ _09503_ vssd1 vssd1 vccd1 vccd1 _09504_ sky130_fd_sc_hd__nor2_1
X_12085_ _04785_ net23 vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__nor2_1
XFILLER_81_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18701_ rbzero.debug_overlay.vplaneY\[0\] vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__buf_2
XFILLER_237_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15913_ _08525_ _08526_ vssd1 vssd1 vccd1 vccd1 _08527_ sky130_fd_sc_hd__or2_1
XFILLER_172_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11036_ _03757_ _03761_ _03763_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__a21bo_1
X_16893_ _07553_ _07837_ vssd1 vssd1 vccd1 vccd1 _09435_ sky130_fd_sc_hd__nand2_1
XFILLER_133_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19681_ rbzero.debug_overlay.playerY\[2\] rbzero.debug_overlay.playerY\[1\] _03032_
+ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__or3_1
XFILLER_237_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15844_ _08109_ _08169_ _08035_ vssd1 vssd1 vccd1 vccd1 _08458_ sky130_fd_sc_hd__a21oi_1
X_18632_ _03736_ rbzero.map_rom.f1 _02356_ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__o21a_1
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15775_ _07517_ _08335_ vssd1 vssd1 vccd1 vccd1 _08389_ sky130_fd_sc_hd__nor2_1
XFILLER_40_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18563_ _02274_ _02191_ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__nor2_1
XFILLER_224_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12987_ _05671_ _05673_ _05674_ _05675_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__a22o_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17514_ _09022_ _08851_ _09373_ _08890_ vssd1 vssd1 vccd1 vccd1 _10051_ sky130_fd_sc_hd__o22ai_1
X_14726_ rbzero.debug_overlay.playerX\[-6\] vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__inv_2
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18494_ _02226_ _02236_ _02240_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__a21oi_2
X_11938_ _04623_ _04647_ _04648_ _04639_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__a22o_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17445_ _09977_ _09981_ _09982_ vssd1 vssd1 vccd1 vccd1 _09983_ sky130_fd_sc_hd__nand3_1
XFILLER_32_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14657_ _03800_ _07300_ _07301_ _07257_ vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__o211a_1
XFILLER_53_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11869_ rbzero.tex_b1\[1\] rbzero.tex_b1\[0\] _03934_ vssd1 vssd1 vccd1 vccd1 _04583_
+ sky130_fd_sc_hd__mux2_1
XFILLER_220_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13608_ _06242_ _06275_ _06277_ _06296_ _06273_ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__o221a_1
XFILLER_177_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17376_ _09828_ _09844_ vssd1 vssd1 vccd1 vccd1 _09914_ sky130_fd_sc_hd__or2_1
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14588_ _07248_ vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__buf_2
XFILLER_201_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16327_ _08798_ _08800_ vssd1 vssd1 vccd1 vccd1 _08938_ sky130_fd_sc_hd__nor2_1
XFILLER_174_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19115_ _09243_ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__buf_4
XFILLER_199_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13539_ _06226_ _06227_ vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__nand2_1
XFILLER_158_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19046_ _02684_ vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__clkbuf_1
X_16258_ _08867_ _08868_ vssd1 vssd1 vccd1 vccd1 _08869_ sky130_fd_sc_hd__xor2_1
XFILLER_220_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15209_ _04933_ _07820_ _07821_ _07822_ vssd1 vssd1 vccd1 vccd1 _07823_ sky130_fd_sc_hd__a31o_1
XFILLER_173_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16189_ _08798_ _08800_ vssd1 vssd1 vccd1 vccd1 _08801_ sky130_fd_sc_hd__xor2_1
XFILLER_142_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19948_ _03114_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__buf_4
XFILLER_228_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19879_ _03110_ vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__clkinv_2
XFILLER_68_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20723_ net93 _00739_ vssd1 vssd1 vccd1 vccd1 rbzero.othery\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20654_ net63 _00670_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20585_ net95 _00601_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21206_ _00255_ _01222_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21137_ _00186_ _01153_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21068_ _00117_ _01084_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12910_ _05350_ _05430_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__nor2_1
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20019_ _03124_ vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__clkinv_2
XFILLER_59_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13890_ _06317_ _06541_ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__or2_1
XFILLER_74_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12841_ _05528_ _05529_ _05444_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__mux2_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15560_ _07467_ _07575_ vssd1 vssd1 vccd1 vccd1 _08174_ sky130_fd_sc_hd__nor2_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12772_ _05454_ _05457_ _05460_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__mux2_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _05602_ _07086_ _07124_ _07177_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_14_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ rbzero.tex_g1\[34\] _03959_ _03916_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__a21o_1
XFILLER_226_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15491_ _08101_ _08103_ _08104_ vssd1 vssd1 vccd1 vccd1 _08105_ sky130_fd_sc_hd__a21o_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _09769_ vssd1 vssd1 vccd1 vccd1 _09770_ sky130_fd_sc_hd__inv_2
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _07105_ _05499_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__nor2_1
XFILLER_159_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11654_ rbzero.color_sky\[2\] rbzero.color_floor\[2\] _04030_ vssd1 vssd1 vccd1 vccd1
+ _04371_ sky130_fd_sc_hd__mux2_1
Xfanout70 net72 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__buf_2
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout81 net83 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__buf_2
X_17161_ _09163_ _07837_ _09700_ vssd1 vssd1 vccd1 vccd1 _09701_ sky130_fd_sc_hd__and3_1
X_10605_ rbzero.tex_g1\[59\] rbzero.tex_g1\[60\] _03519_ vssd1 vssd1 vccd1 vccd1 _03522_
+ sky130_fd_sc_hd__mux2_1
Xfanout92 net98 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__buf_2
XFILLER_196_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14373_ _05408_ _07061_ vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__nor2_1
XFILLER_155_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11585_ _04302_ vssd1 vssd1 vccd1 vccd1 o_rgb[7] sky130_fd_sc_hd__buf_4
XFILLER_200_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16112_ _08723_ vssd1 vssd1 vccd1 vccd1 _08724_ sky130_fd_sc_hd__clkbuf_4
XFILLER_183_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13324_ _06006_ _06011_ _06012_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__o21a_1
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17092_ _09382_ _09496_ _09632_ vssd1 vssd1 vccd1 vccd1 _09633_ sky130_fd_sc_hd__a21oi_1
XFILLER_196_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10536_ _03485_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16043_ _08614_ _08655_ vssd1 vssd1 vccd1 vccd1 _08656_ sky130_fd_sc_hd__xnor2_1
XFILLER_196_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13255_ _05893_ _05943_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10467_ _03449_ vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12206_ o_tex_sclk _04873_ _04874_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__a21oi_1
XFILLER_108_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13186_ _05762_ _05778_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__nor2_1
XFILLER_151_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10398_ _03388_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__clkbuf_4
XFILLER_83_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19802_ _03101_ vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_215_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12137_ _04836_ net29 vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__nor2_1
XFILLER_111_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17994_ _01774_ _01775_ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__and2_1
XFILLER_111_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19733_ _03060_ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__buf_2
X_16945_ _09196_ _09216_ _09486_ vssd1 vssd1 vccd1 vccd1 _09487_ sky130_fd_sc_hd__a21o_1
X_12068_ _04768_ _04519_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__nor2_1
XFILLER_42_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11019_ _03742_ _03743_ _03744_ _03745_ _03746_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__o2111a_1
XFILLER_38_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19664_ rbzero.debug_overlay.playerY\[-3\] _03016_ _03026_ _02978_ vssd1 vssd1 vccd1
+ vccd1 _00981_ sky130_fd_sc_hd__o211a_1
X_16876_ _09416_ _09417_ vssd1 vssd1 vccd1 vccd1 _09418_ sky130_fd_sc_hd__nor2_1
XFILLER_231_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18615_ _03798_ _02348_ _02349_ _02350_ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__a31o_1
XFILLER_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15827_ _08352_ _08416_ _08440_ vssd1 vssd1 vccd1 vccd1 _08441_ sky130_fd_sc_hd__a21oi_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19595_ _02956_ _02972_ _02973_ _02780_ vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__o211a_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15758_ _08365_ _08367_ _08371_ vssd1 vssd1 vccd1 vccd1 _08372_ sky130_fd_sc_hd__o21ai_1
X_18546_ _02277_ _02280_ _02288_ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__nand3_1
XFILLER_244_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14709_ rbzero.wall_tracer.stepDistX\[9\] _07237_ _04931_ vssd1 vssd1 vccd1 vccd1
+ _07329_ sky130_fd_sc_hd__mux2_1
XFILLER_178_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15689_ _08273_ _08302_ vssd1 vssd1 vccd1 vccd1 _08303_ sky130_fd_sc_hd__xnor2_1
XFILLER_166_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18477_ _02223_ _02224_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__or2_1
X_17428_ _08760_ _08917_ vssd1 vssd1 vccd1 vccd1 _09966_ sky130_fd_sc_hd__nor2_1
XFILLER_33_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17359_ _09890_ _09891_ _09889_ vssd1 vssd1 vccd1 vccd1 _09897_ sky130_fd_sc_hd__a21boi_1
XFILLER_174_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20370_ net97 _00403_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.b6 sky130_fd_sc_hd__dfxtp_1
XFILLER_107_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19029_ rbzero.pov.spi_buffer\[61\] rbzero.pov.ready_buffer\[61\] _02673_ vssd1 vssd1
+ vccd1 vccd1 _02676_ sky130_fd_sc_hd__mux2_1
XFILLER_134_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20706_ net99 _00722_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20637_ net55 _00653_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ rbzero.row_render.size\[2\] gpout0.hpos\[2\] _04085_ _04088_ vssd1 vssd1
+ vccd1 vccd1 _04089_ sky130_fd_sc_hd__a211o_1
X_20568_ net137 _00584_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10321_ _03370_ vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20499_ net128 _00515_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13040_ _05607_ _05728_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__or2_1
X_10252_ _03334_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10183_ _03295_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__inv_2
XFILLER_65_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14991_ _07581_ _07582_ vssd1 vssd1 vccd1 vccd1 _07605_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13942_ _06574_ _06628_ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__xnor2_1
X_16730_ _09279_ _09280_ _09281_ _09283_ vssd1 vssd1 vccd1 vccd1 _09284_ sky130_fd_sc_hd__a31o_1
XFILLER_75_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16661_ rbzero.row_render.side _09255_ _09258_ _07343_ vssd1 vssd1 vccd1 vccd1 _00497_
+ sky130_fd_sc_hd__a22o_1
X_13873_ _06505_ _06561_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__nor2_1
XFILLER_234_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15612_ _08225_ _08224_ vssd1 vssd1 vccd1 vccd1 _08226_ sky130_fd_sc_hd__xnor2_2
XFILLER_28_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18400_ rbzero.debug_overlay.vplaneX\[-6\] rbzero.wall_tracer.rayAddendX\[-6\] _02153_
+ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a21o_1
XFILLER_210_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12824_ _05379_ _05389_ _05463_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__mux2_1
XFILLER_62_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16592_ _07843_ _09200_ vssd1 vssd1 vccd1 vccd1 _09201_ sky130_fd_sc_hd__nor2_1
X_19380_ _02860_ vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__clkinv_2
XFILLER_222_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18331_ rbzero.wall_tracer.trackDistY\[3\] _02039_ _02094_ _09888_ vssd1 vssd1 vccd1
+ vccd1 _00580_ sky130_fd_sc_hd__o22a_1
XFILLER_167_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15543_ _08154_ _08156_ vssd1 vssd1 vccd1 vccd1 _08157_ sky130_fd_sc_hd__and2_1
XFILLER_163_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12755_ _05359_ _05410_ _05437_ _05443_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__nor4_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18262_ _02027_ _02029_ _02028_ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__a21boi_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11706_ rbzero.tex_g1\[55\] _03964_ _03965_ _03997_ vssd1 vssd1 vccd1 vccd1 _04422_
+ sky130_fd_sc_hd__a31o_1
XFILLER_202_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15474_ _08082_ _08083_ vssd1 vssd1 vccd1 vccd1 _08088_ sky130_fd_sc_hd__nor2_1
X_12686_ _05249_ _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__xnor2_4
XFILLER_124_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17213_ _09627_ _09629_ vssd1 vssd1 vccd1 vccd1 _09753_ sky130_fd_sc_hd__nor2_1
X_14425_ _07011_ _07059_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__or2_1
X_18193_ _01933_ _01972_ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__xnor2_1
XFILLER_202_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11637_ rbzero.tex_g0\[41\] rbzero.tex_g0\[40\] _04000_ vssd1 vssd1 vccd1 vccd1 _04354_
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17144_ _08086_ vssd1 vssd1 vccd1 vccd1 _09684_ sky130_fd_sc_hd__buf_2
X_14356_ _06985_ _07041_ _07044_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__o21a_1
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11568_ rbzero.debug_overlay.playerY\[1\] _04234_ _04209_ rbzero.debug_overlay.playerY\[-3\]
+ _04285_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__a221o_1
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13307_ _05953_ _05969_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17075_ _09479_ _09477_ vssd1 vssd1 vccd1 vccd1 _09616_ sky130_fd_sc_hd__or2b_1
XFILLER_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10519_ _03476_ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14287_ _06372_ _06399_ _06401_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__or3b_1
XFILLER_13_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11499_ _04203_ _04216_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__nor2_1
XFILLER_226_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16026_ _08627_ _08638_ vssd1 vssd1 vccd1 vccd1 _08639_ sky130_fd_sc_hd__xnor2_2
XFILLER_170_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13238_ _05926_ _05902_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13169_ _05743_ _05754_ _05857_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__a21bo_1
XFILLER_135_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17977_ _01644_ _01627_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__or2b_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19716_ _02727_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__buf_2
X_16928_ _04938_ rbzero.wall_tracer.stepDistX\[9\] vssd1 vssd1 vccd1 vccd1 _09470_
+ sky130_fd_sc_hd__nand2_4
XFILLER_111_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19647_ _03442_ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__buf_4
XFILLER_226_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16859_ _09391_ _09400_ vssd1 vssd1 vccd1 vccd1 _09401_ sky130_fd_sc_hd__nand2_1
XFILLER_81_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19578_ _02956_ _02959_ _02961_ _02780_ vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__o211a_1
XFILLER_20_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18529_ _02250_ _02257_ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__or2_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20422_ net123 _00453_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_140_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20353_ gpout2.clk_div\[0\] _03003_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__nor2_1
XFILLER_134_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20284_ _03257_ vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__clkinv_2
XFILLER_162_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10870_ rbzero.tex_b0\[62\] rbzero.tex_b0\[61\] _03660_ vssd1 vssd1 vccd1 vccd1 _03661_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _03815_ _05085_ _05228_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__a21o_1
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12471_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__nand2_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14210_ _06826_ _06884_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11422_ rbzero.tex_r1\[43\] rbzero.tex_r1\[42\] _03980_ vssd1 vssd1 vccd1 vccd1 _04140_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15190_ _07802_ _07803_ vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14141_ _06814_ _06824_ vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__xor2_1
XFILLER_153_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11353_ rbzero.row_render.size\[7\] _04046_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ _03361_ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__clkbuf_1
X_14072_ _06736_ _06760_ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11284_ rbzero.tex_r0\[31\] _03939_ _03941_ _03942_ vssd1 vssd1 vccd1 vccd1 _04003_
+ sky130_fd_sc_hd__a31o_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17900_ _01651_ _01682_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__xor2_1
X_13023_ _05699_ _05701_ _05709_ _05711_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__a31o_1
XFILLER_156_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10235_ _03325_ vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__clkbuf_1
X_18880_ _02593_ vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__clkbuf_1
XTAP_6730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17831_ _01507_ _01509_ _01508_ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__o21bai_1
XFILLER_121_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17762_ _01533_ _01544_ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__or2_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14974_ _07476_ _07490_ _07587_ vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__a21o_1
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19501_ _02918_ vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__clkbuf_1
X_16713_ _09268_ vssd1 vssd1 vccd1 vccd1 _09269_ sky130_fd_sc_hd__clkbuf_4
XFILLER_235_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13925_ _06610_ _06613_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17693_ _01471_ _01476_ _01477_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__nand3_1
XFILLER_208_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19432_ _02882_ vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__clkbuf_1
XFILLER_228_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13856_ _06543_ _06544_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__or2b_1
X_16644_ _09249_ vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_223_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12807_ _05321_ _05383_ _05429_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__mux2_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19363_ _02859_ vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__clkinv_2
X_16575_ _09182_ _07834_ _09040_ _09183_ _08905_ vssd1 vssd1 vccd1 vccd1 _09184_ sky130_fd_sc_hd__o32ai_2
X_13787_ _06469_ _06474_ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__nand2_1
XFILLER_188_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10999_ rbzero.vga_sync.vsync vssd1 vssd1 vccd1 vccd1 o_vsync sky130_fd_sc_hd__clkinv_4
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18314_ _02075_ _02076_ _02077_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__a21o_1
XFILLER_37_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15526_ _08137_ _08138_ vssd1 vssd1 vccd1 vccd1 _08140_ sky130_fd_sc_hd__nor2_1
X_12738_ _05410_ _05415_ _05426_ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__and3b_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19294_ rbzero.spi_registers.got_new_vshift _02742_ _02740_ _02825_ vssd1 vssd1 vccd1
+ vccd1 _00806_ sky130_fd_sc_hd__a31o_1
XFILLER_188_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18245_ rbzero.wall_tracer.trackDistY\[-9\] _01996_ _02020_ _09302_ vssd1 vssd1 vccd1
+ vccd1 _00568_ sky130_fd_sc_hd__o22a_1
X_15457_ _08056_ _08070_ vssd1 vssd1 vccd1 vccd1 _08071_ sky130_fd_sc_hd__and2b_1
XFILLER_148_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12669_ _05351_ _05335_ _05344_ _05357_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__and4bb_1
XFILLER_15_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14408_ _07092_ _07093_ _07094_ _07095_ _07096_ vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__o41a_1
XFILLER_175_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18176_ _01954_ _01955_ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__xor2_1
XFILLER_198_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15388_ _07981_ _07999_ _08001_ vssd1 vssd1 vccd1 vccd1 _08002_ sky130_fd_sc_hd__a21oi_2
XFILLER_156_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17127_ _09665_ _09666_ vssd1 vssd1 vccd1 vccd1 _09667_ sky130_fd_sc_hd__xnor2_2
X_14339_ _05408_ _06991_ _07006_ _07027_ vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__a31oi_4
XFILLER_144_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17058_ _09596_ _09597_ _09591_ vssd1 vssd1 vccd1 vccd1 _09599_ sky130_fd_sc_hd__a21oi_1
XFILLER_171_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16009_ _08620_ _08621_ vssd1 vssd1 vccd1 vccd1 _08622_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20971_ net71 _00987_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20405_ net119 _00436_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_147_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21385_ net113 _01401_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20336_ _02287_ _02150_ _03268_ _03260_ rbzero.wall_tracer.rayAddendX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__a32o_1
XFILLER_107_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20267_ _03255_ vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__clkinv_2
XTAP_6037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20198_ _03216_ _03219_ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ _04666_ _04673_ _04680_ net17 vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__a22o_1
XFILLER_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13710_ _06395_ _06396_ _06398_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__a21oi_1
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10922_ rbzero.tex_b0\[37\] rbzero.tex_b0\[36\] _03682_ vssd1 vssd1 vccd1 vccd1 _03688_
+ sky130_fd_sc_hd__mux2_1
XFILLER_229_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14690_ _07319_ vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__clkbuf_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13641_ _06222_ _06259_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__xnor2_2
XFILLER_147_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10853_ rbzero.tex_g0\[6\] rbzero.tex_g0\[5\] _03649_ vssd1 vssd1 vccd1 vccd1 _03652_
+ sky130_fd_sc_hd__mux2_1
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _08853_ _08861_ vssd1 vssd1 vccd1 vccd1 _08970_ sky130_fd_sc_hd__or2b_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13572_ _06224_ _06258_ _06256_ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__a21o_1
XFILLER_158_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10784_ _03615_ vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__clkbuf_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15311_ _07908_ _07909_ _07923_ vssd1 vssd1 vccd1 vccd1 _07925_ sky130_fd_sc_hd__and3_1
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12523_ rbzero.wall_tracer.visualWallDist\[-2\] _05190_ rbzero.wall_tracer.rcp_sel\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__a21o_1
XFILLER_34_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ _08885_ _08901_ vssd1 vssd1 vccd1 vccd1 _08902_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18030_ _01801_ _01811_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__xnor2_1
X_15242_ _07852_ _07853_ _07855_ vssd1 vssd1 vccd1 vccd1 _07856_ sky130_fd_sc_hd__nand3_1
XFILLER_173_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12454_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[11\] vssd1
+ vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__nand2_2
XFILLER_200_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11405_ rbzero.tex_r1\[55\] rbzero.tex_r1\[54\] _04119_ vssd1 vssd1 vccd1 vccd1 _04123_
+ sky130_fd_sc_hd__mux2_1
X_15173_ _07785_ _07786_ vssd1 vssd1 vccd1 vccd1 _07787_ sky130_fd_sc_hd__nand2_1
XFILLER_158_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12385_ _05076_ _05077_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__and2_1
XFILLER_197_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14124_ _06774_ _06773_ _06757_ vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__a21o_1
X_11336_ rbzero.row_render.size\[3\] vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__inv_2
X_19981_ _03114_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__buf_4
XFILLER_180_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14055_ _06698_ _06742_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__nor2_1
X_18932_ rbzero.pov.spi_buffer\[15\] rbzero.pov.ready_buffer\[15\] _02618_ vssd1 vssd1
+ vccd1 vccd1 _02625_ sky130_fd_sc_hd__mux2_1
XFILLER_180_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11267_ _03956_ _03967_ _03973_ _03983_ _03985_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__o311a_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13006_ _05691_ _05694_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10218_ _03316_ vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__clkbuf_1
X_18863_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[0\] vssd1
+ vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__or2_1
XTAP_6560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11198_ _03912_ _03913_ _03916_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__mux2_1
XTAP_6571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17814_ _01596_ _01597_ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__xnor2_1
XFILLER_223_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18794_ rbzero.wall_tracer.rayAddendY\[5\] _02515_ _03811_ vssd1 vssd1 vccd1 vccd1
+ _02516_ sky130_fd_sc_hd__mux2_1
XFILLER_208_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17745_ _09166_ _08979_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__nor2_1
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14957_ _07568_ _07570_ _07408_ vssd1 vssd1 vccd1 vccd1 _07571_ sky130_fd_sc_hd__a21o_2
XFILLER_94_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13908_ _06526_ _06596_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17676_ _10100_ _01460_ vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__nand2_1
XFILLER_39_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14888_ _07213_ _07156_ _07346_ vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__a21o_1
XFILLER_90_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19415_ _02873_ vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__clkbuf_1
X_16627_ _09096_ _09098_ _09235_ vssd1 vssd1 vccd1 vccd1 _09236_ sky130_fd_sc_hd__o21ba_1
XFILLER_165_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13839_ _06313_ _06342_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__nor2_1
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19346_ _02857_ vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__clkinv_2
X_16558_ _08595_ _09166_ vssd1 vssd1 vccd1 vccd1 _09167_ sky130_fd_sc_hd__nor2_1
XFILLER_143_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15509_ _04936_ _07733_ vssd1 vssd1 vccd1 vccd1 _08123_ sky130_fd_sc_hd__nor2_2
XFILLER_149_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19277_ rbzero.spi_registers.new_other\[10\] rbzero.spi_registers.spi_buffer\[10\]
+ _02812_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__mux2_1
X_16489_ _09096_ _09098_ vssd1 vssd1 vccd1 vccd1 _09099_ sky130_fd_sc_hd__xor2_4
XFILLER_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18228_ _02003_ _02004_ _01998_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__a21bo_1
XFILLER_248_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18159_ _01840_ _01841_ _01838_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__a21oi_1
XFILLER_144_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21170_ _00219_ _01186_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20121_ _03148_ _03151_ _03149_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__a21boi_1
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20052_ _03128_ vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__clkinv_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20954_ net71 _00970_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20885_ net56 _00901_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12170_ net38 net37 _04875_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__and3_1
X_21368_ _00391_ _01384_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11121_ _03836_ _03839_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__nor2_1
XFILLER_218_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20319_ rbzero.traced_texVinit\[8\] _03260_ _09267_ _09507_ vssd1 vssd1 vccd1 vccd1
+ _01402_ sky130_fd_sc_hd__a22o_1
X_21299_ net133 _01315_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ _03730_ _03779_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__nor2_1
XFILLER_192_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15860_ _07217_ _07221_ _07225_ _07687_ vssd1 vssd1 vccd1 vccd1 _08474_ sky130_fd_sc_hd__or4_2
XTAP_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14811_ _07416_ _07424_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__or2_1
XTAP_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15791_ _08388_ _08403_ vssd1 vssd1 vccd1 vccd1 _08405_ sky130_fd_sc_hd__xnor2_1
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17530_ _10065_ _10066_ vssd1 vssd1 vccd1 vccd1 _10067_ sky130_fd_sc_hd__and2_1
XFILLER_205_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14742_ _07352_ vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__buf_4
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11954_ net16 vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__buf_2
XFILLER_205_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10905_ rbzero.tex_b0\[45\] rbzero.tex_b0\[44\] _03671_ vssd1 vssd1 vccd1 vccd1 _03679_
+ sky130_fd_sc_hd__mux2_1
Xtop_ew_algofoogle_148 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_148/HI o_rgb[8] sky130_fd_sc_hd__conb_1
X_17461_ _09973_ _09997_ _09998_ vssd1 vssd1 vccd1 vccd1 _09999_ sky130_fd_sc_hd__and3_1
XFILLER_189_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14673_ _07310_ vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11885_ rbzero.row_render.side _04593_ _04594_ _04595_ _04597_ vssd1 vssd1 vccd1
+ vccd1 _04598_ sky130_fd_sc_hd__o221a_1
XFILLER_233_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_159 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_159/HI o_rgb[21]
+ sky130_fd_sc_hd__conb_1
XFILLER_232_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19200_ _02727_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__buf_4
X_16412_ _08223_ vssd1 vssd1 vccd1 vccd1 _09022_ sky130_fd_sc_hd__buf_2
X_13624_ _05749_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__clkbuf_4
X_10836_ rbzero.tex_g0\[14\] rbzero.tex_g0\[13\] _03638_ vssd1 vssd1 vccd1 vccd1 _03643_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17392_ _09919_ _09929_ vssd1 vssd1 vccd1 vccd1 _09930_ sky130_fd_sc_hd__nand2_1
XFILLER_164_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19131_ rbzero.othery\[2\] _02723_ _02735_ _02728_ vssd1 vssd1 vccd1 vccd1 _00739_
+ sky130_fd_sc_hd__o211a_1
XFILLER_201_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16343_ _08819_ _08821_ _08817_ vssd1 vssd1 vccd1 vccd1 _08954_ sky130_fd_sc_hd__o21a_1
X_13555_ _06242_ _06243_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__and2_1
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10767_ rbzero.tex_g0\[47\] rbzero.tex_g0\[46\] _03605_ vssd1 vssd1 vccd1 vccd1 _03607_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12506_ _05143_ _05194_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__nand2_1
X_16274_ _08769_ _08777_ _08884_ vssd1 vssd1 vccd1 vccd1 _08885_ sky130_fd_sc_hd__a21o_1
XFILLER_201_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19062_ _02693_ vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__clkbuf_1
XFILLER_200_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13486_ _06166_ _06174_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__or2_1
XFILLER_146_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10698_ _03570_ vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18013_ _01779_ _01794_ vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__xor2_1
XFILLER_201_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15225_ _07663_ _07680_ _07837_ _07838_ vssd1 vssd1 vccd1 vccd1 _07839_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_139_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12437_ _05121_ _05126_ _05127_ _05128_ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__a31o_1
XFILLER_154_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15156_ _07768_ _07769_ vssd1 vssd1 vccd1 vccd1 _07770_ sky130_fd_sc_hd__xor2_1
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12368_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[9\] vssd1
+ vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__nand2_1
XFILLER_126_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14107_ _06777_ _06754_ _06776_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__nand3_1
X_11319_ _03938_ _03940_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__and2_1
XFILLER_236_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15087_ _07699_ _07700_ vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__or2_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19964_ _03119_ vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__clkinv_2
X_12299_ rbzero.wall_tracer.trackDistX\[9\] _04991_ _04992_ rbzero.wall_tracer.trackDistX\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__o22a_1
XFILLER_141_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14038_ _06713_ _06714_ _06725_ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__nand3_1
XFILLER_68_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18915_ rbzero.pov.spi_buffer\[7\] rbzero.pov.ready_buffer\[7\] _02608_ vssd1 vssd1
+ vccd1 vccd1 _02616_ sky130_fd_sc_hd__mux2_1
XTAP_7080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19895_ _03112_ vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__clkinv_2
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18846_ _02510_ rbzero.wall_tracer.rayAddendY\[9\] _02558_ vssd1 vssd1 vccd1 vccd1
+ _02563_ sky130_fd_sc_hd__a21o_1
XTAP_6390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18777_ _02472_ rbzero.debug_overlay.vplaneY\[-3\] vssd1 vssd1 vccd1 vccd1 _02499_
+ sky130_fd_sc_hd__and2_1
X_15989_ _07742_ _07552_ _07550_ _07736_ vssd1 vssd1 vccd1 vccd1 _08602_ sky130_fd_sc_hd__or4_1
XFILLER_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17728_ rbzero.wall_tracer.trackDistX\[6\] _09275_ _01506_ _01512_ vssd1 vssd1 vccd1
+ vccd1 _00559_ sky130_fd_sc_hd__o22a_1
XFILLER_236_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17659_ _01429_ _01443_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20670_ net74 _00686_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_189_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19329_ _02856_ vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__clkinv_2
XFILLER_17_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21222_ _00271_ _01238_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21153_ _00202_ _01169_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20104_ _03138_ _03139_ _03135_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__a21bo_1
XFILLER_132_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21084_ _00133_ _01100_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20035_ _03126_ vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__clkinv_2
XFILLER_219_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20937_ net93 _00953_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.mosi_buffer\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_215_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11670_ _04384_ _04385_ _03968_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__mux2_1
XFILLER_187_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20868_ net54 _00884_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10621_ _03388_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__clkbuf_4
XFILLER_167_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20799_ _00017_ _00815_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13340_ _06028_ _05818_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__nand2_1
XFILLER_126_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10552_ rbzero.tex_r0\[21\] rbzero.tex_r0\[20\] _03490_ vssd1 vssd1 vccd1 vccd1 _03494_
+ sky130_fd_sc_hd__mux2_1
XFILLER_127_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13271_ _05611_ _05959_ _05911_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__o21a_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10483_ rbzero.tex_r0\[54\] rbzero.tex_r0\[53\] _03457_ vssd1 vssd1 vccd1 vccd1 _03458_
+ sky130_fd_sc_hd__mux2_1
X_15010_ _07519_ _07602_ vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__or2_1
XFILLER_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12222_ _04923_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12153_ net32 net31 vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__nor2_1
XFILLER_64_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11104_ gpout0.hpos\[5\] _03782_ _03804_ gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1
+ _03823_ sky130_fd_sc_hd__a31o_1
XFILLER_68_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16961_ _08972_ _09228_ _09502_ vssd1 vssd1 vccd1 vccd1 _09503_ sky130_fd_sc_hd__a21oi_1
XFILLER_133_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12084_ _04779_ _04783_ _04791_ net23 vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__a22o_1
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18700_ _02417_ _02420_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__nand2_1
XFILLER_238_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15912_ _08501_ _08502_ _08524_ vssd1 vssd1 vccd1 vccd1 _08526_ sky130_fd_sc_hd__a21oi_1
XFILLER_172_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11035_ _03736_ _03733_ _03752_ _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__or4_1
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19680_ rbzero.debug_overlay.playerY\[1\] _03008_ _03038_ _02989_ vssd1 vssd1 vccd1
+ vccd1 _00985_ sky130_fd_sc_hd__a211o_1
X_16892_ _07553_ _08485_ vssd1 vssd1 vccd1 vccd1 _09434_ sky130_fd_sc_hd__and2_1
XFILLER_231_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18631_ _02364_ vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15843_ _08112_ _08219_ _08454_ _08456_ vssd1 vssd1 vccd1 vccd1 _08457_ sky130_fd_sc_hd__a22o_2
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18562_ _02301_ _02302_ _02299_ _02300_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__o211ai_2
X_15774_ _08364_ _08387_ vssd1 vssd1 vccd1 vccd1 _08388_ sky130_fd_sc_hd__xnor2_1
X_12986_ _05488_ _05658_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__xnor2_1
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17513_ _09952_ _09972_ vssd1 vssd1 vccd1 vccd1 _10050_ sky130_fd_sc_hd__nand2_1
XFILLER_217_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14725_ rbzero.debug_overlay.playerY\[-6\] vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__inv_2
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18493_ _02223_ _02239_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__xnor2_1
X_11937_ net49 net40 net39 net41 _04618_ _04611_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__mux4_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _09182_ _09463_ _09979_ _09980_ vssd1 vssd1 vccd1 vccd1 _09982_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14656_ _05290_ _03800_ vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__nand2_1
X_11868_ rbzero.tex_b1\[2\] _03903_ _03928_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__a21o_1
XFILLER_205_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13607_ _06239_ _06295_ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__nand2_1
X_10819_ rbzero.tex_g0\[22\] rbzero.tex_g0\[21\] _03627_ vssd1 vssd1 vccd1 vccd1 _03634_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17375_ _09807_ _09822_ _09820_ vssd1 vssd1 vccd1 vccd1 _09913_ sky130_fd_sc_hd__a21o_1
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14587_ _07245_ _07247_ _07250_ _07251_ vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__o211a_1
XFILLER_14_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11799_ _03900_ _04501_ _04505_ _03985_ _04513_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__o311a_1
XFILLER_229_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19114_ rbzero.spi_registers.new_other\[6\] _02725_ vssd1 vssd1 vccd1 vccd1 _02726_
+ sky130_fd_sc_hd__or2_1
X_16326_ _08927_ _08936_ vssd1 vssd1 vccd1 vccd1 _08937_ sky130_fd_sc_hd__xor2_1
XFILLER_192_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13538_ _06212_ _06210_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__or2b_1
XFILLER_185_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19045_ rbzero.pov.spi_buffer\[69\] rbzero.pov.ready_buffer\[69\] _02607_ vssd1 vssd1
+ vccd1 vccd1 _02684_ sky130_fd_sc_hd__mux2_1
X_16257_ _08510_ _08735_ vssd1 vssd1 vccd1 vccd1 _08868_ sky130_fd_sc_hd__nor2_1
X_13469_ _06024_ _06026_ _06065_ _06155_ _06157_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__a32o_1
XFILLER_146_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15208_ _07694_ vssd1 vssd1 vccd1 vccd1 _07822_ sky130_fd_sc_hd__inv_2
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16188_ _07843_ _08645_ _08643_ _08799_ vssd1 vssd1 vccd1 vccd1 _08800_ sky130_fd_sc_hd__o31a_1
XFILLER_126_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15139_ _07750_ _07752_ vssd1 vssd1 vccd1 vccd1 _07753_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19947_ _03117_ vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__clkinv_2
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19878_ _03110_ vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__clkinv_2
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18829_ _02509_ _02428_ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__or2_1
XFILLER_56_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20722_ net101 _00738_ vssd1 vssd1 vccd1 vccd1 rbzero.othery\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_224_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20653_ net62 _00669_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20584_ net95 _00600_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21205_ _00254_ _01221_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21136_ _00185_ _01152_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21067_ _00116_ _01083_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20018_ _03124_ vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__clkinv_2
XFILLER_219_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12840_ _05375_ _05372_ _05448_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__mux2_1
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _05459_ _05445_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__nand2_1
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ _07190_ vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__clkbuf_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ rbzero.tex_g1\[35\] _03939_ _03941_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__and3_1
XFILLER_199_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15490_ _08075_ _08100_ vssd1 vssd1 vccd1 vccd1 _08104_ sky130_fd_sc_hd__nor2_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14441_ _07126_ _07128_ _05527_ vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11653_ _04026_ _04318_ _04336_ _04352_ _04369_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__o32a_1
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout60 net73 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_2
Xfanout71 net72 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10604_ _03521_ vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__clkbuf_1
X_17160_ _07472_ _09428_ vssd1 vssd1 vccd1 vccd1 _09700_ sky130_fd_sc_hd__nor2_1
X_14372_ _07029_ _07060_ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__nand2_1
XFILLER_174_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout82 net83 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout93 net94 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_2
X_11584_ _03826_ _04194_ _04301_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__o21ba_1
XFILLER_167_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16111_ _08722_ vssd1 vssd1 vccd1 vccd1 _08723_ sky130_fd_sc_hd__clkbuf_4
X_13323_ _06001_ _06005_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__or2b_1
XFILLER_127_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10535_ rbzero.tex_r0\[29\] rbzero.tex_r0\[28\] _03479_ vssd1 vssd1 vccd1 vccd1 _03485_
+ sky130_fd_sc_hd__mux2_1
X_17091_ _09493_ _09495_ vssd1 vssd1 vccd1 vccd1 _09632_ sky130_fd_sc_hd__nor2_1
XFILLER_128_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16042_ _08653_ _08654_ vssd1 vssd1 vccd1 vccd1 _08655_ sky130_fd_sc_hd__xor2_1
X_13254_ _05612_ _05567_ _05748_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__and3_1
XFILLER_129_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10466_ rbzero.tex_r0\[62\] rbzero.tex_r0\[61\] _03446_ vssd1 vssd1 vccd1 vccd1 _03449_
+ sky130_fd_sc_hd__mux2_1
XFILLER_237_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12205_ gpout5.clk_div\[1\] net51 net53 net52 _04883_ _04873_ vssd1 vssd1 vccd1 vccd1
+ _04911_ sky130_fd_sc_hd__mux4_1
XFILLER_108_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ _05872_ _05873_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__and2_1
XFILLER_100_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10397_ _03410_ vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__clkbuf_1
X_19801_ _03099_ _04920_ _03100_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__and3b_1
XFILLER_233_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12136_ _04830_ _04834_ _04842_ net29 vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__a22o_1
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17993_ _01772_ _01773_ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__nand2_1
XFILLER_69_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19732_ rbzero.pov.ready_buffer\[30\] _03056_ _03059_ rbzero.debug_overlay.facingY\[-1\]
+ _03065_ vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__o221a_1
X_16944_ _09214_ _09215_ vssd1 vssd1 vccd1 vccd1 _09486_ sky130_fd_sc_hd__nor2_1
X_12067_ net24 net25 vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__nand2_1
XFILLER_133_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11018_ rbzero.map_rom.f1 vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__inv_2
X_19663_ rbzero.pov.ready_buffer\[50\] _02958_ _03007_ _03025_ vssd1 vssd1 vccd1 vccd1
+ _03026_ sky130_fd_sc_hd__a211o_1
XFILLER_226_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16875_ _09413_ _09415_ vssd1 vssd1 vccd1 vccd1 _09417_ sky130_fd_sc_hd__and2_1
XFILLER_38_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18614_ rbzero.debug_overlay.playerX\[1\] _04940_ vssd1 vssd1 vccd1 vccd1 _02350_
+ sky130_fd_sc_hd__and2_1
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15826_ _08413_ _08439_ _08415_ vssd1 vssd1 vccd1 vccd1 _08440_ sky130_fd_sc_hd__o21a_1
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19594_ _07410_ _02960_ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__nand2_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18545_ _02247_ rbzero.wall_tracer.rayAddendX\[6\] vssd1 vssd1 vccd1 vccd1 _02288_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_234_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15757_ _07792_ _07843_ _08369_ _08370_ vssd1 vssd1 vccd1 vccd1 _08371_ sky130_fd_sc_hd__o31a_1
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _05627_ _05582_ _05657_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__or3_2
XFILLER_79_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14708_ _07328_ vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_233_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18476_ rbzero.debug_overlay.vplaneX\[-3\] rbzero.debug_overlay.vplaneX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__and2_1
X_15688_ _08275_ _08301_ vssd1 vssd1 vccd1 vccd1 _08302_ sky130_fd_sc_hd__xnor2_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17427_ _09836_ _09961_ _09962_ _09964_ vssd1 vssd1 vccd1 vccd1 _09965_ sky130_fd_sc_hd__a22o_1
XFILLER_221_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14639_ _04985_ _07246_ _07249_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__o21ai_1
XFILLER_18_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17358_ rbzero.wall_tracer.trackDistX\[4\] rbzero.wall_tracer.stepDistX\[4\] vssd1
+ vssd1 vccd1 vccd1 _09896_ sky130_fd_sc_hd__and2_1
XFILLER_147_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16309_ _07229_ _07234_ _08474_ _07237_ vssd1 vssd1 vccd1 vccd1 _08920_ sky130_fd_sc_hd__o31a_1
XFILLER_88_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17289_ _09718_ _09726_ _09827_ vssd1 vssd1 vccd1 vccd1 _09828_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19028_ _02675_ vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20705_ net99 _00721_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20636_ net54 _00652_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20567_ net137 _00583_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10320_ rbzero.tex_b1\[0\] rbzero.tex_b1\[1\] _03366_ vssd1 vssd1 vccd1 vccd1 _03370_
+ sky130_fd_sc_hd__mux2_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20498_ net127 _00514_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ rbzero.tex_b1\[33\] rbzero.tex_b1\[34\] _03333_ vssd1 vssd1 vccd1 vccd1 _03334_
+ sky130_fd_sc_hd__mux2_1
XFILLER_180_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10182_ gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__buf_2
XFILLER_121_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21119_ _00168_ _01135_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_6967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14990_ _07596_ _07603_ vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13941_ _06573_ _06629_ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__nand2_1
XFILLER_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16660_ _09257_ vssd1 vssd1 vccd1 vccd1 _09258_ sky130_fd_sc_hd__clkbuf_4
X_13872_ _06507_ _06556_ _06560_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__o21a_1
XFILLER_75_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15611_ _07697_ _07579_ vssd1 vssd1 vccd1 vccd1 _08225_ sky130_fd_sc_hd__nand2_1
XFILLER_216_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12823_ _05467_ _05500_ _05511_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__o21ai_1
X_16591_ _07453_ rbzero.wall_tracer.stepDistY\[11\] _07694_ _09199_ vssd1 vssd1 vccd1
+ vccd1 _09200_ sky130_fd_sc_hd__a22oi_4
XFILLER_28_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18330_ _05121_ _02092_ _02093_ _02013_ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__a31o_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15542_ _08062_ _08155_ vssd1 vssd1 vccd1 vccd1 _08156_ sky130_fd_sc_hd__and2b_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12754_ _05439_ _05372_ _05440_ _05441_ _05442_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__a311o_1
XFILLER_131_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18261_ rbzero.wall_tracer.trackDistY\[-6\] rbzero.wall_tracer.stepDistY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__and2_1
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ rbzero.tex_g1\[54\] _04374_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__and2_1
X_15473_ _08086_ _07842_ vssd1 vssd1 vccd1 vccd1 _08087_ sky130_fd_sc_hd__nor2_1
X_12685_ _05305_ _05261_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__nand2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17212_ _09660_ _09751_ vssd1 vssd1 vccd1 vccd1 _09752_ sky130_fd_sc_hd__xnor2_1
XFILLER_230_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14424_ _07111_ _07112_ _07105_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__mux2_1
XFILLER_30_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11636_ rbzero.tex_g0\[43\] rbzero.tex_g0\[42\] _04000_ vssd1 vssd1 vccd1 vccd1 _04353_
+ sky130_fd_sc_hd__mux2_1
X_18192_ _01937_ _01971_ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__xnor2_1
XFILLER_168_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17143_ _09681_ _09682_ vssd1 vssd1 vccd1 vccd1 _09683_ sky130_fd_sc_hd__nand2_1
X_14355_ _05586_ _07042_ _07043_ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__or3_1
XFILLER_156_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11567_ rbzero.debug_overlay.playerY\[-2\] _04245_ _04243_ rbzero.debug_overlay.playerY\[0\]
+ _04284_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__a221o_1
XFILLER_144_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13306_ _05992_ _05994_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__nor2_1
XFILLER_143_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10518_ rbzero.tex_r0\[37\] rbzero.tex_r0\[36\] _03468_ vssd1 vssd1 vccd1 vccd1 _03476_
+ sky130_fd_sc_hd__mux2_1
X_17074_ _09606_ _09614_ vssd1 vssd1 vccd1 vccd1 _09615_ sky130_fd_sc_hd__xnor2_1
X_14286_ _06455_ _06974_ vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__nand2_1
XFILLER_144_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11498_ _04210_ _04215_ gpout0.hpos\[4\] vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__or3b_1
XFILLER_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16025_ _08635_ _08637_ vssd1 vssd1 vccd1 vccd1 _08638_ sky130_fd_sc_hd__nand2_1
X_13237_ _05883_ _05884_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__nor2_1
XFILLER_226_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10449_ rbzero.tex_r1\[3\] rbzero.tex_r1\[4\] _03433_ vssd1 vssd1 vccd1 vccd1 _03438_
+ sky130_fd_sc_hd__mux2_1
XFILLER_100_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13168_ _05753_ _05744_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__or2b_1
XFILLER_170_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12119_ net32 _04824_ _04825_ net29 vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__and4b_1
X_17976_ _01668_ _01681_ _01757_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__a21o_1
X_13099_ _05692_ _05640_ _05679_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__and3_1
XFILLER_242_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19715_ rbzero.pov.ready_buffer\[37\] _03056_ _03059_ rbzero.debug_overlay.facingX\[-5\]
+ _03031_ vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__o221a_1
X_16927_ _09461_ _09468_ vssd1 vssd1 vccd1 vccd1 _09469_ sky130_fd_sc_hd__xnor2_1
XFILLER_211_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19646_ _07427_ _02835_ _03012_ _03013_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__o211a_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16858_ _09398_ _09399_ vssd1 vssd1 vccd1 vccd1 _09400_ sky130_fd_sc_hd__and2_1
XFILLER_226_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15809_ _07616_ _07625_ _07680_ _07847_ vssd1 vssd1 vccd1 vccd1 _08423_ sky130_fd_sc_hd__nor4_2
XFILLER_20_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19577_ _02957_ _02960_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__nand2_1
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16789_ _09332_ _09333_ _09334_ vssd1 vssd1 vccd1 vccd1 _09336_ sky130_fd_sc_hd__a21o_1
XFILLER_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18528_ _02272_ vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__clkbuf_1
XFILLER_178_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18459_ _02188_ _02200_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__nand2_1
XFILLER_146_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20421_ net130 _00452_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20352_ rbzero.wall_tracer.rayAddendY\[-6\] _03260_ _09267_ _03278_ vssd1 vssd1 vccd1
+ vccd1 _01417_ sky130_fd_sc_hd__a22o_1
XFILLER_107_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20283_ _04702_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__buf_4
XFILLER_115_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12470_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__or2_1
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11421_ _03932_ _04136_ _04137_ _04138_ _03923_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__o221a_1
XFILLER_32_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20619_ net84 _00635_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14140_ _06828_ vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__inv_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11352_ _04047_ _04070_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__nor2_1
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10303_ rbzero.tex_b1\[8\] rbzero.tex_b1\[9\] _03355_ vssd1 vssd1 vccd1 vccd1 _03361_
+ sky130_fd_sc_hd__mux2_1
X_14071_ _06435_ _06423_ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__nor2_1
XFILLER_152_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11283_ rbzero.tex_r0\[30\] _04001_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__and2_1
XFILLER_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ _05612_ _05710_ _05708_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__and3_1
XFILLER_112_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10234_ rbzero.tex_b1\[41\] rbzero.tex_b1\[42\] _03322_ vssd1 vssd1 vccd1 vccd1 _03325_
+ sky130_fd_sc_hd__mux2_1
XFILLER_106_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17830_ rbzero.wall_tracer.trackDistX\[7\] rbzero.wall_tracer.stepDistX\[7\] vssd1
+ vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__nand2_1
XFILLER_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17761_ _01533_ _01544_ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__nand2_1
XFILLER_43_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14973_ _07532_ _07586_ vssd1 vssd1 vccd1 vccd1 _07587_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19500_ rbzero.pov.spi_buffer\[46\] rbzero.pov.spi_buffer\[47\] _02910_ vssd1 vssd1
+ vccd1 vccd1 _02918_ sky130_fd_sc_hd__mux2_1
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16712_ _03728_ _03809_ vssd1 vssd1 vccd1 vccd1 _09268_ sky130_fd_sc_hd__or2_1
XFILLER_235_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13924_ _06516_ _06611_ _06612_ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__a21bo_1
X_17692_ _01474_ _01475_ _10111_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__a21o_1
XFILLER_48_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19431_ rbzero.pov.spi_buffer\[13\] rbzero.pov.spi_buffer\[14\] _02877_ vssd1 vssd1
+ vccd1 vccd1 _02882_ sky130_fd_sc_hd__mux2_1
X_16643_ _09247_ _04107_ _09248_ vssd1 vssd1 vccd1 vccd1 _09249_ sky130_fd_sc_hd__and3_1
XFILLER_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13855_ _06479_ _06539_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__xor2_1
XFILLER_228_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ _05494_ _05420_ _05429_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__mux2_1
X_19362_ _02859_ vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__clkinv_2
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16574_ _08771_ _08788_ vssd1 vssd1 vccd1 vccd1 _09183_ sky130_fd_sc_hd__nand2_1
XFILLER_76_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13786_ _06469_ _06474_ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__or2_1
X_10998_ _03727_ vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18313_ _02078_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__inv_2
XFILLER_128_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15525_ _08137_ _08138_ vssd1 vssd1 vccd1 vccd1 _08139_ sky130_fd_sc_hd__xor2_2
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12737_ _05416_ _05419_ _05421_ _05424_ _05425_ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__o2111a_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19293_ _02831_ vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18244_ _01997_ _02018_ _02019_ _02013_ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a31o_1
XFILLER_188_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15456_ _08066_ _08068_ _08069_ vssd1 vssd1 vccd1 vccd1 _08070_ sky130_fd_sc_hd__o21ai_1
X_12668_ _05346_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__inv_2
XFILLER_124_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14407_ _07075_ _05408_ vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__nand2_1
XFILLER_89_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18175_ _08536_ _08633_ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__nand2_1
X_11619_ _03899_ _04322_ _04327_ _03985_ _04335_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__o311a_1
X_15387_ _07636_ _08000_ vssd1 vssd1 vccd1 vccd1 _08001_ sky130_fd_sc_hd__or2_1
XFILLER_106_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12599_ _05188_ _05287_ _03790_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__a21o_1
XFILLER_237_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17126_ _07505_ _07506_ _09389_ vssd1 vssd1 vccd1 vccd1 _09666_ sky130_fd_sc_hd__and3_2
XFILLER_15_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14338_ _07007_ _07026_ vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__and2_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17057_ _09591_ _09596_ _09597_ vssd1 vssd1 vccd1 vccd1 _09598_ sky130_fd_sc_hd__and3_1
X_14269_ _06851_ _06957_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__xnor2_1
XFILLER_217_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16008_ _07751_ _07712_ vssd1 vssd1 vccd1 vccd1 _08621_ sky130_fd_sc_hd__nor2_1
XFILLER_135_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17959_ _07631_ _08634_ _01739_ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__o21ai_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20970_ net71 _00986_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_226_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19629_ rbzero.debug_overlay.playerX\[4\] _02995_ vssd1 vssd1 vccd1 vccd1 _03000_
+ sky130_fd_sc_hd__and2b_1
XFILLER_241_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20404_ net119 _00435_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_147_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21384_ net112 _01400_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20335_ _02147_ _02149_ _02148_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__a21bo_1
XFILLER_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20266_ _03255_ vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__clkinv_2
XTAP_6016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20197_ _03217_ _03218_ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__and2b_1
XFILLER_0_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _04664_ net18 _04674_ _04676_ _04679_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__a32o_1
XFILLER_245_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10921_ _03687_ vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13640_ _06324_ _06328_ _06316_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__a21o_1
X_10852_ _03651_ vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _06222_ _06259_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__nor2_2
X_10783_ rbzero.tex_g0\[39\] rbzero.tex_g0\[38\] _03605_ vssd1 vssd1 vccd1 vccd1 _03615_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15310_ _07908_ _07909_ _07923_ vssd1 vssd1 vccd1 vccd1 _07924_ sky130_fd_sc_hd__a21oi_1
XFILLER_164_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12522_ _03789_ _05210_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__nand2_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _08892_ _08900_ vssd1 vssd1 vccd1 vccd1 _08901_ sky130_fd_sc_hd__xor2_2
XFILLER_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15241_ _07683_ _07714_ _07854_ vssd1 vssd1 vccd1 vccd1 _07855_ sky130_fd_sc_hd__a21o_1
XFILLER_36_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12453_ _05142_ vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11404_ _04120_ _04121_ _03909_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__mux2_1
XFILLER_201_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15172_ _07774_ _07778_ vssd1 vssd1 vccd1 vccd1 _07786_ sky130_fd_sc_hd__or2b_1
XFILLER_166_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12384_ _05030_ _05031_ _05075_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__nand3_1
XFILLER_181_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14123_ _06774_ _06757_ _06773_ vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__nand3_1
X_11335_ rbzero.row_render.size\[4\] vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__inv_2
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19980_ _03120_ vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__clkinv_2
XFILLER_153_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18931_ _02624_ vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__clkbuf_1
X_14054_ _06310_ _06542_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__nor2_1
XFILLER_10_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11266_ _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__buf_6
XFILLER_107_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13005_ _05692_ _05618_ _05693_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__o21ai_1
X_10217_ rbzero.tex_b1\[49\] rbzero.tex_b1\[50\] _03311_ vssd1 vssd1 vccd1 vccd1 _03316_
+ sky130_fd_sc_hd__mux2_1
XFILLER_239_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18862_ rbzero.spi_registers.spi_counter\[6\] rbzero.spi_registers.spi_counter\[5\]
+ rbzero.spi_registers.spi_counter\[4\] vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__or3_1
XTAP_6550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11197_ _03915_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__buf_6
XFILLER_84_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17813_ _01470_ _01484_ _01482_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__a21o_1
XTAP_6572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18793_ _03729_ _02504_ _02514_ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__a21o_1
XFILLER_223_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17744_ _09684_ _08852_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__nor2_1
XTAP_5882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14956_ _07334_ _05247_ _07569_ vssd1 vssd1 vccd1 vccd1 _07570_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13907_ _06313_ _06389_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__nor2_1
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17675_ _08923_ _09470_ _08241_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__a21oi_1
XFILLER_235_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14887_ _04937_ _07491_ _07495_ _07500_ vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__a31oi_4
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19414_ rbzero.pov.spi_buffer\[5\] rbzero.pov.spi_buffer\[6\] _02866_ vssd1 vssd1
+ vccd1 vccd1 _02873_ sky130_fd_sc_hd__mux2_1
X_16626_ _08955_ _09095_ vssd1 vssd1 vccd1 vccd1 _09235_ sky130_fd_sc_hd__and2b_1
X_13838_ _06310_ _06330_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__or2_1
XFILLER_63_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19345_ _02857_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__clkinv_2
XFILLER_204_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16557_ _07936_ vssd1 vssd1 vccd1 vccd1 _09166_ sky130_fd_sc_hd__buf_2
XFILLER_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13769_ _06441_ _06439_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__xor2_1
XFILLER_204_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15508_ _07467_ _07485_ vssd1 vssd1 vccd1 vccd1 _08122_ sky130_fd_sc_hd__nor2_1
XFILLER_188_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19276_ _02822_ vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16488_ _08710_ _08827_ _08958_ _09097_ _08957_ vssd1 vssd1 vccd1 vccd1 _09098_ sky130_fd_sc_hd__a32oi_4
XFILLER_104_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18227_ _01998_ _02003_ _02004_ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__nand3b_1
X_15439_ _08042_ _08044_ _08052_ vssd1 vssd1 vccd1 vccd1 _08053_ sky130_fd_sc_hd__o21ai_1
XFILLER_164_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18158_ _01872_ _01881_ _01879_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a21bo_1
XFILLER_157_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17109_ _09631_ _09633_ vssd1 vssd1 vccd1 vccd1 _09649_ sky130_fd_sc_hd__or2_1
XFILLER_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18089_ _01868_ _01869_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__nor2_1
XFILLER_144_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20120_ rbzero.traced_texa\[-8\] rbzero.texV\[-8\] vssd1 vssd1 vccd1 vccd1 _03154_
+ sky130_fd_sc_hd__and2_1
XFILLER_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20051_ _03128_ vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__clkinv_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20953_ net91 _00969_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ net58 _00900_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21367_ _00390_ _01383_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_218_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11120_ rbzero.texV\[5\] _03837_ _03838_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__a21boi_1
XFILLER_162_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20318_ _02197_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__clkbuf_4
XFILLER_150_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21298_ net114 _01314_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11051_ _03731_ _03778_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__or2_1
XFILLER_89_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20249_ _03253_ vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__clkinv_2
XFILLER_103_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _07423_ vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__buf_2
XTAP_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15790_ _08388_ _08403_ vssd1 vssd1 vccd1 vccd1 _08404_ sky130_fd_sc_hd__nor2_1
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14741_ _07350_ _07353_ _07354_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__a21o_2
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11953_ _04622_ _04642_ _04662_ _04663_ vssd1 vssd1 vccd1 vccd1 o_gpout[1] sky130_fd_sc_hd__o31a_4
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17460_ _09994_ _09995_ _09996_ vssd1 vssd1 vccd1 vccd1 _09998_ sky130_fd_sc_hd__a21o_1
XFILLER_205_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10904_ _03678_ vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__clkbuf_1
XFILLER_229_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14672_ rbzero.wall_tracer.stepDistX\[-9\] _07157_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _07310_ sky130_fd_sc_hd__mux2_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_149 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_149/HI o_rgb[9] sky130_fd_sc_hd__conb_1
X_11884_ _03288_ _04596_ rbzero.row_render.wall\[0\] _04592_ vssd1 vssd1 vccd1 vccd1
+ _04597_ sky130_fd_sc_hd__a211o_1
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16411_ _08223_ _07598_ _09020_ vssd1 vssd1 vccd1 vccd1 _09021_ sky130_fd_sc_hd__or3_1
XFILLER_233_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13623_ _06311_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__inv_2
X_17391_ _09927_ _09928_ vssd1 vssd1 vccd1 vccd1 _09929_ sky130_fd_sc_hd__and2_1
X_10835_ _03642_ vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19130_ rbzero.spi_registers.new_other\[2\] _02725_ vssd1 vssd1 vccd1 vccd1 _02735_
+ sky130_fd_sc_hd__or2_1
X_16342_ _08846_ _08952_ vssd1 vssd1 vccd1 vccd1 _08953_ sky130_fd_sc_hd__xnor2_1
X_13554_ _06238_ _06201_ _06241_ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__or3_1
XFILLER_158_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10766_ _03606_ vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12505_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[11\] vssd1
+ vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__or2_1
X_19061_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.spi_buffer\[1\]
+ _02690_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__mux2_1
X_16273_ _08770_ _08776_ vssd1 vssd1 vccd1 vccd1 _08884_ sky130_fd_sc_hd__and2b_1
XFILLER_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13485_ _06167_ _06173_ vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__and2_1
XFILLER_173_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10697_ rbzero.tex_g1\[15\] rbzero.tex_g1\[16\] _03563_ vssd1 vssd1 vccd1 vccd1 _03570_
+ sky130_fd_sc_hd__mux2_1
XFILLER_160_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18012_ _01792_ _01793_ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__nor2_1
XFILLER_200_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15224_ rbzero.debug_overlay.playerX\[-9\] _04937_ _07643_ vssd1 vssd1 vccd1 vccd1
+ _07838_ sky130_fd_sc_hd__a21o_4
XFILLER_145_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12436_ rbzero.debug_overlay.playerY\[2\] _04940_ vssd1 vssd1 vccd1 vccd1 _05128_
+ sky130_fd_sc_hd__and2_1
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15155_ _07742_ _07468_ vssd1 vssd1 vccd1 vccd1 _07769_ sky130_fd_sc_hd__nor2_1
X_12367_ _05059_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__inv_2
XFILLER_99_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14106_ _06733_ _06781_ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__xor2_2
XFILLER_153_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ rbzero.floor_leak\[5\] _03896_ _03984_ rbzero.floor_leak\[4\] vssd1 vssd1
+ vccd1 vccd1 _04037_ sky130_fd_sc_hd__o22a_1
X_12298_ rbzero.wall_tracer.trackDistY\[8\] vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__inv_2
X_15086_ _07470_ _07685_ _07696_ _07471_ vssd1 vssd1 vccd1 vccd1 _07700_ sky130_fd_sc_hd__o22a_1
X_19963_ _03119_ vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__clkinv_2
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14037_ _06713_ _06714_ _06725_ vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__a21o_1
X_11249_ _03916_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__buf_4
X_18914_ _02615_ vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__clkbuf_1
XTAP_7070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19894_ _03112_ vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__clkinv_2
XTAP_7092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18845_ rbzero.wall_tracer.rayAddendY\[9\] _03812_ _09269_ _02560_ _02562_ vssd1
+ vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__o221a_1
XTAP_6380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18776_ _02472_ rbzero.debug_overlay.vplaneY\[-3\] vssd1 vssd1 vccd1 vccd1 _02498_
+ sky130_fd_sc_hd__nor2_1
XFILLER_227_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15988_ _08598_ _08600_ vssd1 vssd1 vccd1 vccd1 _08601_ sky130_fd_sc_hd__xnor2_2
XTAP_5690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17727_ _09303_ _01510_ _01511_ _09282_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__a31o_1
X_14939_ _07550_ vssd1 vssd1 vccd1 vccd1 _07553_ sky130_fd_sc_hd__clkinv_4
XFILLER_247_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17658_ _01441_ _01442_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__nor2_1
XFILLER_247_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16609_ _09069_ _09071_ vssd1 vssd1 vccd1 vccd1 _09218_ sky130_fd_sc_hd__and2_1
XFILLER_211_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17589_ _10122_ _10123_ _10125_ vssd1 vssd1 vccd1 vccd1 _10126_ sky130_fd_sc_hd__nand3_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19328_ _02856_ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__clkinv_2
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19259_ rbzero.spi_registers.new_other\[0\] rbzero.spi_registers.spi_buffer\[0\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__mux2_1
XFILLER_108_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21221_ _00270_ _01237_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21152_ _00201_ _01168_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20103_ _03135_ _03138_ _03139_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__nand3b_1
XFILLER_99_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21083_ _00132_ _01099_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20034_ _03126_ vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__clkinv_2
XFILLER_101_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ net70 _00952_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[73\] sky130_fd_sc_hd__dfxtp_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20867_ net79 _00883_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10620_ _03529_ vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20798_ net86 _00814_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10551_ _03493_ vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13270_ _05627_ _05657_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__or2_4
X_10482_ _03445_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__clkbuf_4
XFILLER_211_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12221_ o_vsync rbzero.wall_tracer.state\[7\] _04920_ vssd1 vssd1 vccd1 vccd1 _04923_
+ sky130_fd_sc_hd__and3_1
XFILLER_120_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12152_ net31 net32 vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__and2b_1
XFILLER_163_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11103_ gpout0.vpos\[2\] gpout0.vpos\[1\] gpout0.vpos\[0\] _03821_ gpout0.vpos\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__o41a_1
XFILLER_46_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16960_ _09226_ _09227_ vssd1 vssd1 vccd1 vccd1 _09502_ sky130_fd_sc_hd__nor2_1
X_12083_ _04773_ net24 _04784_ _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__a31o_1
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15911_ _08501_ _08502_ _08524_ vssd1 vssd1 vccd1 vccd1 _08525_ sky130_fd_sc_hd__and3_1
X_11034_ rbzero.map_rom.d6 _03744_ rbzero.map_rom.i_row\[4\] _03758_ vssd1 vssd1 vccd1
+ vccd1 _03762_ sky130_fd_sc_hd__or4_1
XFILLER_77_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16891_ _09431_ _09432_ vssd1 vssd1 vccd1 vccd1 _09433_ sky130_fd_sc_hd__xnor2_2
XFILLER_238_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18630_ rbzero.map_rom.f1 _02363_ _09274_ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__mux2_1
X_15842_ _08112_ _08455_ vssd1 vssd1 vccd1 vccd1 _08456_ sky130_fd_sc_hd__xnor2_1
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18561_ _02299_ _02300_ _02301_ _02302_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a211o_1
XFILLER_246_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15773_ _08373_ _08372_ vssd1 vssd1 vccd1 vccd1 _08387_ sky130_fd_sc_hd__and2b_1
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12985_ _05604_ _05659_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__nor2_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17512_ _09954_ _09971_ vssd1 vssd1 vccd1 vccd1 _10049_ sky130_fd_sc_hd__or2_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _07337_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__buf_4
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18492_ _02237_ _02238_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__nor2_1
X_11936_ net42 net44 net43 _04116_ net9 _04618_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__mux4_1
XFILLER_220_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17443_ _07858_ _09463_ _09979_ _09980_ vssd1 vssd1 vccd1 vccd1 _09981_ sky130_fd_sc_hd__or4bb_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14655_ rbzero.wall_tracer.trackDistX\[8\] rbzero.wall_tracer.trackDistY\[8\] _05025_
+ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__mux2_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ rbzero.tex_b1\[3\] _03859_ _03901_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__and3_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13606_ _06231_ _06294_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17374_ _09782_ _09911_ vssd1 vssd1 vccd1 vccd1 _09912_ sky130_fd_sc_hd__xnor2_2
XFILLER_159_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10818_ _03633_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14586_ _03819_ vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__buf_2
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11798_ _03924_ _04508_ _04512_ _03950_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__a211o_1
X_19113_ rbzero.spi_registers.got_new_other _02724_ vssd1 vssd1 vccd1 vccd1 _02725_
+ sky130_fd_sc_hd__nand2_2
X_16325_ _08933_ _08935_ vssd1 vssd1 vccd1 vccd1 _08936_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13537_ _06209_ _06181_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__or2b_1
XFILLER_53_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10749_ rbzero.tex_g0\[55\] rbzero.tex_g0\[54\] _03593_ vssd1 vssd1 vccd1 vccd1 _03597_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19044_ _02683_ vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__clkbuf_1
X_16256_ _08865_ _08866_ vssd1 vssd1 vccd1 vccd1 _08867_ sky130_fd_sc_hd__nand2_1
X_13468_ _06024_ _06156_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15207_ _07217_ _07221_ _07687_ vssd1 vssd1 vccd1 vccd1 _07821_ sky130_fd_sc_hd__or3_1
XFILLER_127_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12419_ _05065_ _05066_ _05067_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__a21bo_2
X_16187_ _08641_ _08642_ vssd1 vssd1 vccd1 vccd1 _08799_ sky130_fd_sc_hd__nand2_1
XFILLER_86_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13399_ _06070_ _06082_ _06087_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__a21bo_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15138_ _07469_ _07751_ vssd1 vssd1 vccd1 vccd1 _07752_ sky130_fd_sc_hd__nor2_1
XFILLER_153_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15069_ _07666_ _07682_ vssd1 vssd1 vccd1 vccd1 _07683_ sky130_fd_sc_hd__xor2_1
XFILLER_141_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19946_ _03117_ vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__clkinv_2
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19877_ _03110_ vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__clkinv_2
XFILLER_60_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18828_ _02510_ _02428_ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__nand2_1
XFILLER_228_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18759_ _02464_ _02468_ _02481_ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__nor3_1
XFILLER_83_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20721_ net93 _00737_ vssd1 vssd1 vccd1 vccd1 rbzero.othery\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20652_ net62 _00668_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20583_ net95 _00599_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21204_ _00253_ _01220_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21135_ _00184_ _01151_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21066_ _00115_ _01082_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20017_ _03124_ vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__clkinv_2
XFILLER_98_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12770_ _05458_ _05452_ _05428_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__or3b_2
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ rbzero.tex_g1\[33\] rbzero.tex_g1\[32\] _03980_ vssd1 vssd1 vccd1 vccd1 _04437_
+ sky130_fd_sc_hd__mux2_1
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20919_ net68 _00935_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[56\] sky130_fd_sc_hd__dfxtp_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14440_ _05517_ _07127_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__or2_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _03985_ _04360_ _04368_ _03896_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__a31o_1
XFILLER_74_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout61 net73 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_2
XFILLER_168_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10603_ rbzero.tex_g1\[60\] rbzero.tex_g1\[61\] _03519_ vssd1 vssd1 vccd1 vccd1 _03521_
+ sky130_fd_sc_hd__mux2_1
Xfanout72 net73 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__buf_2
X_14371_ _07016_ _07059_ _05586_ vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__mux2_1
Xfanout83 net98 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_2
XFILLER_161_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout94 net95 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_2
X_11583_ _04116_ _04115_ _04300_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__or3_1
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16110_ _05290_ _08629_ _04938_ vssd1 vssd1 vccd1 vccd1 _08722_ sky130_fd_sc_hd__or3_1
XFILLER_168_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13322_ _06009_ _06010_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__xor2_1
XFILLER_122_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17090_ _09526_ _09630_ vssd1 vssd1 vccd1 vccd1 _09631_ sky130_fd_sc_hd__xnor2_1
XFILLER_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10534_ _03484_ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16041_ _08496_ _08498_ vssd1 vssd1 vccd1 vccd1 _08654_ sky130_fd_sc_hd__and2_1
XFILLER_202_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13253_ _05671_ _05610_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__nor2_1
X_10465_ _03448_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_237_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12204_ _04871_ net35 _04902_ _04906_ _04909_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__a311o_1
XFILLER_108_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13184_ _05843_ _05844_ _05871_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__or3_1
XFILLER_135_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10396_ rbzero.tex_r1\[28\] rbzero.tex_r1\[29\] _03400_ vssd1 vssd1 vccd1 vccd1 _03410_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19800_ gpout0.vpos\[6\] _04104_ _03094_ gpout0.vpos\[7\] vssd1 vssd1 vccd1 vccd1
+ _03100_ sky130_fd_sc_hd__a31o_1
X_12135_ _04825_ net30 _04835_ _04841_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__a31o_1
XFILLER_237_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17992_ _01772_ _01773_ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__or2_1
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16943_ _09460_ _09484_ vssd1 vssd1 vccd1 vccd1 _09485_ sky130_fd_sc_hd__xnor2_1
XFILLER_238_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19731_ rbzero.pov.ready_buffer\[29\] _03056_ _03059_ rbzero.debug_overlay.facingY\[-2\]
+ _03065_ vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__o221a_1
XFILLER_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12066_ net26 _04772_ _04773_ net23 vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__and4b_1
XFILLER_111_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11017_ rbzero.map_rom.f4 rbzero.map_rom.d6 rbzero.map_rom.c6 rbzero.map_rom.f3 vssd1
+ vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__o22a_1
X_16874_ _09413_ _09415_ vssd1 vssd1 vccd1 vccd1 _09416_ sky130_fd_sc_hd__nor2_1
X_19662_ _07534_ _02958_ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__nor2_1
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15825_ _08383_ _08417_ _08386_ _08438_ vssd1 vssd1 vccd1 vccd1 _08439_ sky130_fd_sc_hd__or4b_1
X_18613_ rbzero.map_rom.f4 _02347_ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__nand2_1
XFILLER_168_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19593_ rbzero.pov.ready_buffer\[64\] _07413_ _02962_ vssd1 vssd1 vccd1 vccd1 _02972_
+ sky130_fd_sc_hd__mux2_1
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15756_ _07517_ _08335_ _08368_ vssd1 vssd1 vccd1 vccd1 _08370_ sky130_fd_sc_hd__or3_1
XFILLER_80_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18544_ _09257_ vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__clkbuf_4
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12968_ _05488_ _05471_ _05474_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__and3_2
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14707_ rbzero.wall_tracer.stepDistX\[8\] _07234_ _04931_ vssd1 vssd1 vccd1 vccd1
+ _07328_ sky130_fd_sc_hd__mux2_1
XFILLER_221_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18475_ rbzero.debug_overlay.vplaneX\[-3\] rbzero.debug_overlay.vplaneX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__nor2_1
X_11919_ net12 vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__inv_2
X_15687_ _08274_ _07971_ vssd1 vssd1 vccd1 vccd1 _08301_ sky130_fd_sc_hd__nor2_1
XFILLER_127_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12899_ _05586_ _05547_ _05587_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__a21o_1
XFILLER_209_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _07553_ _09963_ vssd1 vssd1 vccd1 vccd1 _09964_ sky130_fd_sc_hd__nand2_1
X_14638_ _04941_ _07254_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__nor2_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17357_ rbzero.wall_tracer.trackDistX\[4\] rbzero.wall_tracer.stepDistX\[4\] vssd1
+ vssd1 vccd1 vccd1 _09895_ sky130_fd_sc_hd__nor2_1
X_14569_ _05440_ _07007_ _07069_ _07236_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__a31o_2
XFILLER_158_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16308_ _07229_ _07234_ _07237_ _08474_ vssd1 vssd1 vccd1 vccd1 _08919_ sky130_fd_sc_hd__nor4_2
XFILLER_179_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17288_ _09719_ _09725_ vssd1 vssd1 vccd1 vccd1 _09827_ sky130_fd_sc_hd__and2b_1
XFILLER_174_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19027_ rbzero.pov.spi_buffer\[60\] rbzero.pov.ready_buffer\[60\] _02673_ vssd1 vssd1
+ vccd1 vccd1 _02675_ sky130_fd_sc_hd__mux2_1
X_16239_ _08849_ vssd1 vssd1 vccd1 vccd1 _08850_ sky130_fd_sc_hd__buf_2
XFILLER_174_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19929_ _03116_ vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__clkinv_2
XFILLER_102_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20704_ net87 _00720_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20635_ net55 _00651_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20566_ net137 _00582_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20497_ net127 _00513_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10250_ _03299_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10181_ _03293_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__buf_2
XTAP_6924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21118_ _00167_ _01134_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_6957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13940_ _06574_ _06628_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__nand2_1
X_21049_ _00098_ _01065_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13871_ _06557_ _06559_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__or2b_1
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15610_ _08223_ _07971_ vssd1 vssd1 vccd1 vccd1 _08224_ sky130_fd_sc_hd__nor2_2
XFILLER_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12822_ _05360_ _05504_ _05510_ _05481_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__o22a_1
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16590_ _07240_ _09198_ _08919_ _07337_ vssd1 vssd1 vccd1 vccd1 _09199_ sky130_fd_sc_hd__a31o_1
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15541_ _07552_ _08059_ vssd1 vssd1 vccd1 vccd1 _08155_ sky130_fd_sc_hd__nor2_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12753_ _05298_ _05300_ _05307_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__a21boi_1
XFILLER_43_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18260_ rbzero.wall_tracer.trackDistY\[-6\] rbzero.wall_tracer.stepDistY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__nor2_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _04418_ _04419_ _03958_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__mux2_1
XFILLER_231_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15472_ _08085_ vssd1 vssd1 vccd1 vccd1 _08086_ sky130_fd_sc_hd__clkbuf_4
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12684_ _05369_ _05372_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__or2_1
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _09748_ _09750_ vssd1 vssd1 vccd1 vccd1 _09751_ sky130_fd_sc_hd__xor2_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14423_ _07002_ _07018_ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__or2_1
XFILLER_187_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18191_ _01964_ _01970_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__xnor2_1
XFILLER_202_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11635_ _03900_ _04343_ _04351_ _03954_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__o211a_1
XFILLER_30_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17142_ _07617_ _07621_ _07709_ _09166_ vssd1 vssd1 vccd1 vccd1 _09682_ sky130_fd_sc_hd__or4_1
X_14354_ _05432_ _07001_ vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__and2_1
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11566_ gpout0.vpos\[5\] gpout0.vpos\[4\] _04246_ vssd1 vssd1 vccd1 vccd1 _04284_
+ sky130_fd_sc_hd__or3_1
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13305_ _05983_ _05989_ _05991_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__nor3_1
X_17073_ _09612_ _09613_ vssd1 vssd1 vccd1 vccd1 _09614_ sky130_fd_sc_hd__and2b_1
XFILLER_196_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10517_ _03475_ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__clkbuf_1
X_14285_ _06571_ _06973_ _06567_ _06569_ vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__a211o_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11497_ _04198_ _04197_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__or2_1
XFILLER_157_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16024_ _04929_ _07698_ _08633_ _08636_ _07697_ vssd1 vssd1 vccd1 vccd1 _08637_ sky130_fd_sc_hd__a32o_1
XFILLER_157_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13236_ _05906_ _05924_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__nand2_1
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10448_ _03437_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13167_ _05756_ _05855_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10379_ _03401_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__clkbuf_1
X_12118_ net28 vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__buf_2
XFILLER_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17975_ _01678_ _01680_ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__nor2_1
X_13098_ _05692_ _05641_ _05679_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a21oi_1
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19714_ rbzero.pov.ready_buffer\[36\] _03056_ _03059_ rbzero.debug_overlay.facingX\[-6\]
+ _03031_ vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__o221a_1
XFILLER_66_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16926_ _09463_ _09467_ vssd1 vssd1 vccd1 vccd1 _09468_ sky130_fd_sc_hd__nor2_1
X_12049_ _04750_ _04754_ _04757_ _04720_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__a22o_1
XFILLER_120_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19645_ rbzero.pov.ready_buffer\[45\] _02835_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__nand2_1
XFILLER_77_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16857_ _09396_ _09397_ vssd1 vssd1 vccd1 vccd1 _09399_ sky130_fd_sc_hd__nand2_1
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15808_ _08419_ _08421_ vssd1 vssd1 vccd1 vccd1 _08422_ sky130_fd_sc_hd__and2_1
XFILLER_168_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16788_ _09332_ _09333_ _09334_ vssd1 vssd1 vccd1 vccd1 _09335_ sky130_fd_sc_hd__nand3_1
X_19576_ _02955_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__clkbuf_4
XFILLER_241_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15739_ _08351_ _08352_ vssd1 vssd1 vccd1 vccd1 _08353_ sky130_fd_sc_hd__nor2_1
X_18527_ rbzero.wall_tracer.rayAddendX\[4\] _02271_ _03812_ vssd1 vssd1 vccd1 vccd1
+ _02272_ sky130_fd_sc_hd__mux2_1
XFILLER_209_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18458_ _02203_ _02206_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17409_ _09914_ _09846_ _09946_ vssd1 vssd1 vccd1 vccd1 _09947_ sky130_fd_sc_hd__a21o_1
XFILLER_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18389_ rbzero.debug_overlay.vplaneX\[-5\] rbzero.wall_tracer.rayAddendX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__nor2_1
XFILLER_92_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20420_ net123 _00451_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_144_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20351_ _02380_ _03277_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20282_ _03256_ vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__clkinv_2
XFILLER_192_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11420_ rbzero.tex_r1\[47\] _03939_ _03941_ _04014_ vssd1 vssd1 vccd1 vccd1 _04138_
+ sky130_fd_sc_hd__a31o_1
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20618_ net84 _00634_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_240_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11351_ rbzero.row_render.size\[8\] rbzero.row_render.size\[7\] _04046_ vssd1 vssd1
+ vccd1 vccd1 _04070_ sky130_fd_sc_hd__nor3_1
XFILLER_125_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20549_ net124 _00565_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10302_ _03360_ vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__clkbuf_1
X_14070_ _06724_ _06723_ _06716_ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__a21o_1
XFILLER_180_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ _04000_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__buf_4
XFILLER_180_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13021_ _05703_ _05704_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__nand2_1
XFILLER_69_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10233_ _03324_ vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17760_ _01542_ _01543_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__and2_1
X_14972_ _07584_ _07585_ vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__and2b_1
XFILLER_120_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13923_ _06471_ _06470_ _06320_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__or3b_1
XFILLER_169_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16711_ rbzero.traced_texa\[11\] _09266_ _09267_ rbzero.wall_tracer.visualWallDist\[11\]
+ vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__a22o_1
XFILLER_48_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17691_ _10111_ _01474_ _01475_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__nand3_1
XFILLER_235_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16642_ _04591_ _04085_ vssd1 vssd1 vccd1 vccd1 _09248_ sky130_fd_sc_hd__or2_1
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19430_ _02881_ vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__clkbuf_1
X_13854_ _05861_ _06542_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__or2_1
XFILLER_90_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12805_ _05325_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__clkinv_2
X_16573_ _07858_ vssd1 vssd1 vccd1 vccd1 _09182_ sky130_fd_sc_hd__clkbuf_4
X_19361_ _02859_ vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__clkinv_2
X_13785_ _06470_ _06471_ _06473_ _06468_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10997_ rbzero.tex_b0\[1\] rbzero.tex_b0\[0\] _03445_ vssd1 vssd1 vccd1 vccd1 _03727_
+ sky130_fd_sc_hd__mux2_1
X_18312_ _02075_ _02076_ _02077_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__and3_1
X_15524_ _07260_ _07408_ _04935_ _07384_ vssd1 vssd1 vccd1 vccd1 _08138_ sky130_fd_sc_hd__or4_2
XFILLER_71_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12736_ _05361_ _05363_ _05382_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__or3_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19292_ rbzero.spi_registers.new_vshift\[5\] rbzero.spi_registers.spi_buffer\[5\]
+ _02825_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__mux2_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18243_ _02015_ _02016_ _02017_ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a21o_1
XFILLER_148_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15455_ _08058_ _08065_ vssd1 vssd1 vccd1 vccd1 _08069_ sky130_fd_sc_hd__or2_1
XFILLER_128_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12667_ _05310_ _05322_ _05350_ _05355_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__and4_1
XFILLER_19_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14406_ _06990_ _06987_ _07031_ _05568_ vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__a31o_1
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18174_ _07670_ _09389_ vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__nand2_1
XFILLER_15_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11618_ _03921_ _04330_ _04334_ _03950_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__a211o_1
X_15386_ _07622_ _07635_ vssd1 vssd1 vccd1 vccd1 _08000_ sky130_fd_sc_hd__and2_1
XFILLER_128_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12598_ rbzero.wall_tracer.visualWallDist\[5\] _05190_ vssd1 vssd1 vccd1 vccd1 _05287_
+ sky130_fd_sc_hd__nand2_1
XFILLER_50_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17125_ _09663_ _09664_ vssd1 vssd1 vccd1 vccd1 _09665_ sky130_fd_sc_hd__nand2_1
XFILLER_237_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14337_ _07023_ _07025_ _05531_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__mux2_1
XFILLER_128_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11549_ _04262_ _04266_ gpout0.vpos\[5\] _04106_ vssd1 vssd1 vccd1 vccd1 _04267_
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17056_ _09592_ _09594_ _09595_ vssd1 vssd1 vccd1 vccd1 _09597_ sky130_fd_sc_hd__a21o_1
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14268_ _06875_ _06874_ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__nor2_1
XFILLER_125_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16007_ _08463_ _08617_ _08618_ _08619_ vssd1 vssd1 vccd1 vccd1 _08620_ sky130_fd_sc_hd__a22o_1
X_13219_ _05800_ _05799_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__and2b_1
XFILLER_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14199_ _05668_ _06176_ _06387_ _06861_ vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__a31o_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _07631_ _08634_ _01739_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__or3_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16909_ _09450_ vssd1 vssd1 vccd1 vccd1 _09451_ sky130_fd_sc_hd__buf_2
XFILLER_211_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17889_ _10095_ _08671_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__nor2_1
XFILLER_66_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19628_ _02955_ _02998_ rbzero.debug_overlay.playerX\[4\] vssd1 vssd1 vccd1 vccd1
+ _02999_ sky130_fd_sc_hd__o21ai_1
XFILLER_199_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19559_ _02948_ vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20403_ net121 _00434_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
X_21383_ net112 _01399_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20334_ _02287_ _02148_ _03267_ _03260_ rbzero.wall_tracer.rayAddendX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__a32o_1
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20265_ _03255_ vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__clkinv_2
XTAP_6006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20196_ rbzero.traced_texa\[4\] rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1 _03218_
+ sky130_fd_sc_hd__nand2_1
XFILLER_49_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10920_ rbzero.tex_b0\[38\] rbzero.tex_b0\[37\] _03682_ vssd1 vssd1 vccd1 vccd1 _03687_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10851_ rbzero.tex_g0\[7\] rbzero.tex_g0\[6\] _03649_ vssd1 vssd1 vccd1 vccd1 _03651_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _06224_ _06258_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__xor2_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10782_ _03614_ vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__clkbuf_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _05205_ _05209_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__xnor2_2
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15240_ _07666_ _07682_ vssd1 vssd1 vccd1 vccd1 _07854_ sky130_fd_sc_hd__nor2_1
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ _05141_ rbzero.map_rom.i_row\[4\] _05028_ vssd1 vssd1 vccd1 vccd1 _05142_
+ sky130_fd_sc_hd__mux2_1
XFILLER_199_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11403_ rbzero.tex_r1\[51\] rbzero.tex_r1\[50\] _04119_ vssd1 vssd1 vccd1 vccd1 _04121_
+ sky130_fd_sc_hd__mux2_1
X_15171_ _07777_ _07775_ vssd1 vssd1 vccd1 vccd1 _07785_ sky130_fd_sc_hd__or2b_1
XFILLER_138_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12383_ _05031_ _05075_ _05030_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__a21o_1
XFILLER_165_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14122_ _06809_ _06810_ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__nor2_1
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11334_ rbzero.row_render.size\[5\] vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__inv_2
XFILLER_158_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14053_ _06313_ _06542_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__nor2_1
XFILLER_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18930_ rbzero.pov.spi_buffer\[14\] rbzero.pov.ready_buffer\[14\] _02618_ vssd1 vssd1
+ vccd1 vccd1 _02624_ sky130_fd_sc_hd__mux2_1
XFILLER_153_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11265_ _03872_ _03894_ _03952_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__or3_2
XFILLER_180_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13004_ _05608_ _05611_ _05537_ _05635_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__or4_1
XFILLER_49_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10216_ _03315_ vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__clkbuf_1
X_18861_ _02575_ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__clkbuf_2
XTAP_6540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11196_ _03914_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__buf_4
XFILLER_239_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17812_ _01583_ _01595_ vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__xnor2_1
XTAP_6573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18792_ _03818_ _02512_ _02513_ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__and3_1
XFILLER_239_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17743_ _01451_ _01468_ _01526_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__a21o_1
XTAP_5883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14955_ _07341_ _05095_ _07336_ vssd1 vssd1 vccd1 vccd1 _07569_ sky130_fd_sc_hd__o21a_1
XFILLER_212_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13906_ _06266_ _06423_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__nor2_1
X_17674_ _08241_ _09462_ _01458_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__o21a_1
X_14886_ _07496_ _07499_ _07466_ vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__a21oi_2
XFILLER_78_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19413_ _02872_ vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__clkbuf_1
XFILLER_223_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16625_ _09232_ _09233_ vssd1 vssd1 vccd1 vccd1 _09234_ sky130_fd_sc_hd__or2b_2
X_13837_ _06310_ _06342_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__or2_1
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16556_ _09163_ _08893_ _09028_ _09164_ vssd1 vssd1 vccd1 vccd1 _09165_ sky130_fd_sc_hd__a31o_1
XFILLER_189_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19344_ _02857_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__clkinv_2
X_13768_ _06434_ _06443_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12719_ _05407_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__buf_2
X_15507_ _08117_ _08120_ _08118_ vssd1 vssd1 vccd1 vccd1 _08121_ sky130_fd_sc_hd__a21o_1
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16487_ _08840_ _08825_ vssd1 vssd1 vccd1 vccd1 _09097_ sky130_fd_sc_hd__nand2_1
XFILLER_143_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19275_ rbzero.spi_registers.new_other\[9\] rbzero.spi_registers.spi_buffer\[9\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__mux2_1
X_13699_ _06176_ _06387_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__nand2_2
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18226_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.stepDistY\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__nand2_1
X_15438_ _08050_ _08051_ vssd1 vssd1 vccd1 vccd1 _08052_ sky130_fd_sc_hd__or2b_1
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18157_ _01934_ _01936_ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__xnor2_1
X_15369_ _07606_ _07608_ _07609_ vssd1 vssd1 vccd1 vccd1 _07983_ sky130_fd_sc_hd__a21oi_1
XFILLER_156_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17108_ rbzero.wall_tracer.trackDistX\[1\] _09301_ _09641_ _09648_ vssd1 vssd1 vccd1
+ vccd1 _00554_ sky130_fd_sc_hd__o22a_1
X_18088_ _01865_ _01867_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__and2_1
XFILLER_85_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17039_ _09578_ _09579_ vssd1 vssd1 vccd1 vccd1 _09580_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20050_ _03128_ vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__clkinv_2
XFILLER_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20952_ net116 _00968_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_242_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20883_ net58 _00899_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21366_ _00389_ _01382_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20317_ rbzero.traced_texVinit\[7\] _09266_ _09237_ _09261_ vssd1 vssd1 vccd1 vccd1
+ _01401_ sky130_fd_sc_hd__a22o_1
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21297_ net134 _01313_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11050_ _03756_ _03764_ _03777_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__nor3_2
XFILLER_157_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20248_ _03253_ vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__clkinv_2
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20179_ _03199_ _03200_ _03201_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__a21o_1
XFILLER_118_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14740_ _04927_ rbzero.wall_tracer.stepDistX\[-4\] vssd1 vssd1 vccd1 vccd1 _07354_
+ sky130_fd_sc_hd__nor2_1
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ _04658_ o_rgb[15] _04652_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__or3b_1
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10903_ rbzero.tex_b0\[46\] rbzero.tex_b0\[45\] _03671_ vssd1 vssd1 vccd1 vccd1 _03678_
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14671_ _07309_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__clkbuf_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ rbzero.row_render.wall\[1\] vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__inv_2
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16410_ _09017_ _09019_ vssd1 vssd1 vccd1 vccd1 _09020_ sky130_fd_sc_hd__nand2_1
XFILLER_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13622_ _05434_ _06306_ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__nor2_1
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17390_ _09925_ _09926_ vssd1 vssd1 vccd1 vccd1 _09928_ sky130_fd_sc_hd__nand2_1
XFILLER_189_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10834_ rbzero.tex_g0\[15\] rbzero.tex_g0\[14\] _03638_ vssd1 vssd1 vccd1 vccd1 _03642_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16341_ _08949_ _08951_ vssd1 vssd1 vccd1 vccd1 _08952_ sky130_fd_sc_hd__xor2_1
XFILLER_213_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13553_ _06238_ _06201_ _06241_ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__o21ai_2
XFILLER_160_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10765_ rbzero.tex_g0\[48\] rbzero.tex_g0\[47\] _03605_ vssd1 vssd1 vccd1 vccd1 _03606_
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12504_ _05187_ _05192_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__nand2_1
X_19060_ _02692_ vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__clkbuf_1
X_16272_ _08754_ _08762_ _08882_ vssd1 vssd1 vccd1 vccd1 _08883_ sky130_fd_sc_hd__a21o_1
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13484_ _06168_ _06172_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__nand2_1
XFILLER_146_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10696_ _03569_ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18011_ _01789_ _01791_ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__and2_1
X_15223_ _04929_ _07832_ _07651_ _07833_ vssd1 vssd1 vccd1 vccd1 _07837_ sky130_fd_sc_hd__a31o_2
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12435_ _05124_ _05125_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__nand2_1
XFILLER_126_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15154_ _07766_ _07767_ vssd1 vssd1 vccd1 vccd1 _07768_ sky130_fd_sc_hd__and2b_1
X_12366_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[10\] vssd1
+ vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__xor2_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14105_ _06789_ _06793_ vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__or2_1
XFILLER_154_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11317_ rbzero.floor_leak\[3\] _03949_ _03984_ rbzero.floor_leak\[4\] _04035_ vssd1
+ vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__a221o_1
X_15085_ _07685_ _07696_ _07697_ _07698_ vssd1 vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__and4bb_1
X_19962_ _03119_ vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__clkinv_2
X_12297_ rbzero.wall_tracer.trackDistY\[9\] vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__inv_2
XFILLER_153_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14036_ _06716_ _06723_ _06724_ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__a21bo_1
XFILLER_113_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18913_ rbzero.pov.spi_buffer\[6\] rbzero.pov.ready_buffer\[6\] _02608_ vssd1 vssd1
+ vccd1 vccd1 _02615_ sky130_fd_sc_hd__mux2_1
XTAP_7060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11248_ _03958_ _03960_ _03963_ _03966_ _03924_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__o221a_1
XTAP_7071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19893_ _03112_ vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__clkinv_2
XTAP_7082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18844_ _02548_ _02552_ _02561_ _03818_ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__a211o_1
XTAP_6370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11179_ _03868_ _03894_ _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__nor3_4
XTAP_6381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18775_ rbzero.wall_tracer.rayAddendY\[4\] _03812_ _02490_ _02497_ vssd1 vssd1 vccd1
+ vccd1 _00621_ sky130_fd_sc_hd__o22a_1
X_15987_ _08599_ _07598_ vssd1 vssd1 vccd1 vccd1 _08600_ sky130_fd_sc_hd__nor2_1
XTAP_5680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17726_ _01507_ _01508_ _01509_ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__o21ai_1
X_14938_ _07542_ vssd1 vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__buf_2
XFILLER_242_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17657_ _01438_ _01440_ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__and2_1
XFILLER_223_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14869_ _04927_ rbzero.wall_tracer.stepDistX\[-7\] vssd1 vssd1 vccd1 vccd1 _07483_
+ sky130_fd_sc_hd__nor2_2
XFILLER_223_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16608_ _09196_ _09216_ vssd1 vssd1 vccd1 vccd1 _09217_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17588_ _09985_ _09986_ _09993_ _10124_ vssd1 vssd1 vccd1 vccd1 _10125_ sky130_fd_sc_hd__o31ai_1
XFILLER_189_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19327_ _02855_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__buf_4
X_16539_ _09142_ _09147_ vssd1 vssd1 vccd1 vccd1 _09148_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19258_ _02812_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__clkbuf_4
XFILLER_104_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18209_ _01911_ _01915_ _01987_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__or3_1
XFILLER_176_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19189_ rbzero.color_floor\[5\] _02763_ _02772_ vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__a21o_1
XFILLER_191_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21220_ _00269_ _01236_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21151_ _00200_ _01167_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20102_ rbzero.traced_texa\[-11\] rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1 _03139_
+ sky130_fd_sc_hd__nand2_1
X_21082_ _00131_ _01098_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20033_ _03126_ vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__clkinv_2
XFILLER_150_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20935_ net69 _00951_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[72\] sky130_fd_sc_hd__dfxtp_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20866_ net79 _00882_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20797_ net86 _00813_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10550_ rbzero.tex_r0\[22\] rbzero.tex_r0\[21\] _03490_ vssd1 vssd1 vccd1 vccd1 _03493_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10481_ _03456_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12220_ _04922_ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12151_ _04836_ net29 _04851_ _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__a31o_1
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21349_ _00372_ _01365_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11102_ gpout0.vpos\[5\] gpout0.vpos\[4\] gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1
+ _03821_ sky130_fd_sc_hd__or3_2
XFILLER_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12082_ _04785_ _04786_ _04788_ _04789_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__o211a_1
XFILLER_81_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15910_ _08503_ _08523_ vssd1 vssd1 vccd1 vccd1 _08524_ sky130_fd_sc_hd__xnor2_1
X_11033_ _03735_ _03743_ rbzero.map_rom.c6 rbzero.map_rom.f1 _03760_ vssd1 vssd1 vccd1
+ vccd1 _03761_ sky130_fd_sc_hd__o221a_1
XFILLER_133_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16890_ _07598_ _09166_ vssd1 vssd1 vccd1 vccd1 _09432_ sky130_fd_sc_hd__nor2_1
XFILLER_172_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15841_ _08167_ _08219_ vssd1 vssd1 vccd1 vccd1 _08455_ sky130_fd_sc_hd__nor2_1
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18560_ rbzero.wall_tracer.rayAddendX\[6\] rbzero.wall_tracer.rayAddendX\[5\] rbzero.wall_tracer.rayAddendX\[4\]
+ rbzero.wall_tracer.rayAddendX\[3\] _02274_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__o41a_1
XFILLER_224_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15772_ _08377_ _08385_ vssd1 vssd1 vccd1 vccd1 _08386_ sky130_fd_sc_hd__xnor2_1
X_12984_ _05672_ _05624_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__nor2_1
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17511_ _09941_ _09942_ _09944_ vssd1 vssd1 vccd1 vccd1 _10048_ sky130_fd_sc_hd__o21ai_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14723_ _07336_ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__buf_4
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11935_ o_tex_oeb0 _04643_ _04644_ net47 _04645_ vssd1 vssd1 vccd1 vccd1 _04646_
+ sky130_fd_sc_hd__a221o_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18491_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.debug_overlay.vplaneX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__nor2_1
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17442_ _08771_ _09607_ _09611_ _08046_ vssd1 vssd1 vccd1 vccd1 _09980_ sky130_fd_sc_hd__a22o_1
XFILLER_221_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14654_ _03800_ _07298_ _07299_ _07257_ vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__o211a_1
XFILLER_45_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11866_ _04578_ _04579_ _03908_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__mux2_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13605_ _05645_ _05701_ _06270_ _06293_ _05703_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__a32o_1
XFILLER_92_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10817_ rbzero.tex_g0\[23\] rbzero.tex_g0\[22\] _03627_ vssd1 vssd1 vccd1 vccd1 _03633_
+ sky130_fd_sc_hd__mux2_1
X_17373_ _09909_ _09910_ vssd1 vssd1 vccd1 vccd1 _09911_ sky130_fd_sc_hd__nor2_1
XFILLER_232_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14585_ rbzero.wall_tracer.visualWallDist\[-12\] _07249_ vssd1 vssd1 vccd1 vccd1
+ _07250_ sky130_fd_sc_hd__or2_1
XFILLER_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11797_ _03957_ _04509_ _04510_ _04511_ _03946_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__o221a_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19112_ _02721_ vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__clkbuf_4
X_16324_ _08796_ _08797_ _08934_ vssd1 vssd1 vccd1 vccd1 _08935_ sky130_fd_sc_hd__a21oi_1
X_13536_ _06178_ _06216_ vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__and2_1
X_10748_ _03596_ vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_229_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16255_ _08592_ _08732_ _08536_ _08507_ vssd1 vssd1 vccd1 vccd1 _08866_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_201_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19043_ rbzero.pov.spi_buffer\[68\] rbzero.pov.ready_buffer\[68\] _02673_ vssd1 vssd1
+ vccd1 vccd1 _02683_ sky130_fd_sc_hd__mux2_1
XFILLER_173_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13467_ _06026_ _06065_ _06023_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__a21oi_1
XFILLER_220_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10679_ _03560_ vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__clkbuf_1
X_15206_ _07689_ _07690_ _07819_ vssd1 vssd1 vccd1 vccd1 _07820_ sky130_fd_sc_hd__a21o_1
XFILLER_145_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12418_ _05102_ _05106_ _05110_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__or3b_1
XFILLER_86_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16186_ _08796_ _08797_ vssd1 vssd1 vccd1 vccd1 _08798_ sky130_fd_sc_hd__xnor2_1
X_13398_ _06085_ _06086_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__nand2_1
XFILLER_154_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15137_ _07416_ vssd1 vssd1 vccd1 vccd1 _07751_ sky130_fd_sc_hd__clkbuf_4
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12349_ rbzero.debug_overlay.facingY\[-7\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__and2_1
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15068_ _07677_ _07679_ _07681_ vssd1 vssd1 vccd1 vccd1 _07682_ sky130_fd_sc_hd__a21boi_1
XFILLER_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19945_ _03117_ vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__clkinv_2
XFILLER_218_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14019_ _06696_ _06703_ _06705_ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__and3_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19876_ _03110_ vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__clkinv_2
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18827_ _02544_ _02545_ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__xnor2_1
XFILLER_56_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18758_ _02464_ _02468_ _02481_ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__o21a_1
XFILLER_209_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17709_ _10161_ _01493_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__xnor2_1
XFILLER_209_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18689_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__nand2_1
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20720_ net93 _00736_ vssd1 vssd1 vccd1 vccd1 rbzero.otherx\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20651_ net62 _00667_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20582_ net93 _00598_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21203_ _00252_ _01219_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21134_ _00183_ _01150_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21065_ _00114_ _01081_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_235_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20016_ _03124_ vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__clkinv_2
XFILLER_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _04434_ _04435_ _03997_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__mux2_1
XFILLER_226_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20918_ net68 _00934_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11651_ _03921_ _04363_ _04367_ _03899_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__a211o_1
XFILLER_230_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20849_ _00067_ _00865_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10602_ _03520_ vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__clkbuf_1
Xfanout62 net64 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__buf_2
X_14370_ _07058_ vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__inv_2
XFILLER_126_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11582_ _03293_ _03296_ _03807_ _03826_ _04299_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__o311a_1
Xfanout73 net1 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_4
Xfanout84 net89 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__buf_2
XFILLER_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout95 net98 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__buf_2
X_13321_ _05607_ _06007_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__or2_1
XFILLER_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10533_ rbzero.tex_r0\[30\] rbzero.tex_r0\[29\] _03479_ vssd1 vssd1 vccd1 vccd1 _03484_
+ sky130_fd_sc_hd__mux2_1
XFILLER_210_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ _08626_ _08652_ vssd1 vssd1 vccd1 vccd1 _08653_ sky130_fd_sc_hd__xnor2_1
XFILLER_182_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13252_ _05618_ _05745_ _05629_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10464_ rbzero.tex_r0\[63\] rbzero.tex_r0\[62\] _03446_ vssd1 vssd1 vccd1 vccd1 _03448_
+ sky130_fd_sc_hd__mux2_1
XFILLER_237_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12203_ _04873_ _04883_ _04908_ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__nor3_1
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13183_ _05843_ _05844_ _05871_ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__o21ai_1
X_10395_ _03409_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12134_ _04836_ _04837_ _04839_ _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__o211a_1
X_17991_ _07760_ _08725_ _01659_ _01657_ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__o31a_1
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19730_ rbzero.pov.ready_buffer\[28\] _03061_ _03063_ rbzero.debug_overlay.facingY\[-3\]
+ _03066_ vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__a221o_1
X_16942_ _09481_ _09483_ vssd1 vssd1 vccd1 vccd1 _09484_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12065_ net22 vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__buf_2
XFILLER_145_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11016_ rbzero.map_rom.a6 vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__inv_2
X_19661_ rbzero.debug_overlay.playerY\[-4\] _03016_ _03024_ _02978_ vssd1 vssd1 vccd1
+ vccd1 _00980_ sky130_fd_sc_hd__o211a_1
XFILLER_238_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16873_ _09141_ _09148_ _09414_ vssd1 vssd1 vccd1 vccd1 _09415_ sky130_fd_sc_hd__a21oi_1
XFILLER_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18612_ rbzero.map_rom.f4 _02347_ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__or2_1
X_15824_ _08435_ _08436_ _08410_ _08437_ vssd1 vssd1 vccd1 vccd1 _08438_ sky130_fd_sc_hd__and4b_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19592_ _02956_ _02970_ _02971_ _02780_ vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__o211a_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ rbzero.wall_tracer.rayAddendX\[5\] _02158_ _02280_ _02281_ _02286_ vssd1
+ vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__a221o_1
X_15755_ _07517_ _08335_ _08368_ vssd1 vssd1 vccd1 vccd1 _08369_ sky130_fd_sc_hd__o21a_1
X_12967_ _05654_ _05655_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__xor2_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14706_ _07327_ vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__clkbuf_1
X_11918_ gpout0.hpos\[2\] _04080_ _04628_ _04101_ net9 _04625_ vssd1 vssd1 vccd1 vccd1
+ _04629_ sky130_fd_sc_hd__mux4_1
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18474_ _02218_ _02219_ _02220_ _02204_ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__a22o_1
XFILLER_248_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15686_ _08292_ _08299_ vssd1 vssd1 vccd1 vccd1 _08300_ sky130_fd_sc_hd__xnor2_1
XFILLER_166_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12898_ _05586_ _05571_ _05405_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__o21ai_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17425_ _08478_ _08928_ vssd1 vssd1 vccd1 vccd1 _09963_ sky130_fd_sc_hd__nand2_1
X_14637_ _07245_ _07286_ _07287_ _07251_ vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__o211a_1
X_11849_ _04561_ _04562_ _03915_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__mux2_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ _07213_ vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__inv_2
X_17356_ rbzero.wall_tracer.trackDistX\[3\] _09301_ _09888_ _09894_ vssd1 vssd1 vccd1
+ vccd1 _00556_ sky130_fd_sc_hd__o22a_1
XFILLER_147_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16307_ _08629_ rbzero.wall_tracer.stepDistY\[9\] vssd1 vssd1 vccd1 vccd1 _08918_
+ sky130_fd_sc_hd__nand2_1
XFILLER_186_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13519_ _05866_ _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__xor2_1
XFILLER_105_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17287_ _09710_ _09711_ _09713_ vssd1 vssd1 vccd1 vccd1 _09826_ sky130_fd_sc_hd__o21ai_1
XFILLER_179_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14499_ _07181_ vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19026_ _02674_ vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__clkbuf_1
X_16238_ _08629_ _04939_ rbzero.wall_tracer.visualWallDist\[9\] vssd1 vssd1 vccd1
+ vccd1 _08849_ sky130_fd_sc_hd__or3b_1
XFILLER_174_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16169_ _08629_ rbzero.wall_tracer.stepDistY\[8\] vssd1 vssd1 vccd1 vccd1 _08781_
+ sky130_fd_sc_hd__nand2_1
XFILLER_177_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19928_ _03116_ vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__clkinv_2
XFILLER_229_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19859_ _02862_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__buf_4
XFILLER_112_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20703_ net87 _00719_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20634_ net55 _00650_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20565_ net136 _00581_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20496_ net127 _00512_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10180_ gpout0.hpos\[8\] vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__clkbuf_4
XTAP_6914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21117_ _00166_ _01133_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_6958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21048_ _00097_ _01064_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13870_ _06547_ _06552_ _06558_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__a21bo_1
XFILLER_189_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12821_ _05507_ _05509_ _05478_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__mux2_1
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15540_ _08153_ _08064_ vssd1 vssd1 vccd1 vccd1 _08154_ sky130_fd_sc_hd__xnor2_1
X_12752_ _05402_ _05329_ _05335_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__and3_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11703_ rbzero.tex_g1\[51\] rbzero.tex_g1\[50\] _04378_ vssd1 vssd1 vccd1 vccd1 _04419_
+ sky130_fd_sc_hd__mux2_1
X_15471_ _07439_ _07440_ vssd1 vssd1 vccd1 vccd1 _08085_ sky130_fd_sc_hd__and2_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12683_ _05370_ _05371_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__xor2_4
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _09566_ _09626_ _09749_ vssd1 vssd1 vccd1 vccd1 _09750_ sky130_fd_sc_hd__a21oi_1
X_14422_ _07015_ _07021_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__or2b_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _03921_ _04346_ _04350_ _03950_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__a211o_1
X_18190_ _01968_ _01969_ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17141_ rbzero.wall_tracer.visualWallDist\[4\] _03796_ _08123_ _09680_ vssd1 vssd1
+ vccd1 vccd1 _09681_ sky130_fd_sc_hd__a31o_1
X_14353_ _06981_ _07017_ vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__and2_1
XFILLER_50_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11565_ rbzero.debug_overlay.playerY\[2\] _04235_ _04282_ rbzero.debug_overlay.playerY\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__a22o_1
XFILLER_156_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13304_ _05951_ _05972_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17072_ _09609_ _09611_ _09476_ _09608_ vssd1 vssd1 vccd1 vccd1 _09613_ sky130_fd_sc_hd__a211o_1
X_10516_ rbzero.tex_r0\[38\] rbzero.tex_r0\[37\] _03468_ vssd1 vssd1 vccd1 vccd1 _03475_
+ sky130_fd_sc_hd__mux2_1
X_14284_ _06630_ _06690_ _06970_ _06972_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__a31o_1
X_11496_ _04213_ _04207_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__and2_2
XFILLER_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16023_ _08485_ vssd1 vssd1 vccd1 vccd1 _08636_ sky130_fd_sc_hd__buf_2
X_13235_ _05907_ _05922_ _05923_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__a21oi_1
XFILLER_143_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10447_ rbzero.tex_r1\[4\] rbzero.tex_r1\[5\] _03433_ vssd1 vssd1 vccd1 vccd1 _03437_
+ sky130_fd_sc_hd__mux2_1
XFILLER_237_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13166_ _05845_ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__xnor2_1
XFILLER_237_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10378_ rbzero.tex_r1\[37\] rbzero.tex_r1\[38\] _03400_ vssd1 vssd1 vccd1 vccd1 _03401_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12117_ _04820_ o_rgb[7] _04823_ net31 vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__a211o_1
XFILLER_112_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17974_ _01754_ _01755_ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__xor2_1
X_13097_ _05685_ _05785_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__nor2_1
XFILLER_78_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19713_ rbzero.pov.ready_buffer\[35\] _03056_ _03059_ rbzero.debug_overlay.facingX\[-7\]
+ _03031_ vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__o221a_1
X_16925_ _09465_ _09466_ vssd1 vssd1 vccd1 vccd1 _09467_ sky130_fd_sc_hd__nand2_2
X_12048_ net53 _04748_ _04755_ net51 _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__a221o_1
XFILLER_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19644_ net40 _02954_ _02721_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__o21a_2
X_16856_ _09396_ _09397_ vssd1 vssd1 vccd1 vccd1 _09398_ sky130_fd_sc_hd__or2_1
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15807_ _07521_ _08136_ _08395_ _08420_ vssd1 vssd1 vccd1 vccd1 _08421_ sky130_fd_sc_hd__a22o_1
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19575_ _02957_ rbzero.pov.ready_buffer\[59\] _02958_ vssd1 vssd1 vccd1 vccd1 _02959_
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16787_ _09325_ _09327_ _09326_ vssd1 vssd1 vccd1 vccd1 _09334_ sky130_fd_sc_hd__o21bai_1
XFILLER_4_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13999_ _06628_ _06687_ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__nor2_1
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18526_ _02258_ _02259_ _02268_ _02270_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__o22ai_1
X_15738_ _08283_ _08312_ vssd1 vssd1 vccd1 vccd1 _08352_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18457_ _02204_ _02205_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__nand2_1
XFILLER_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15669_ _08282_ _08155_ vssd1 vssd1 vccd1 vccd1 _08283_ sky130_fd_sc_hd__and2b_1
XFILLER_221_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17408_ _09944_ _09945_ vssd1 vssd1 vccd1 vccd1 _09946_ sky130_fd_sc_hd__nand2_1
XFILLER_53_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18388_ _02142_ vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17339_ _09788_ _09877_ vssd1 vssd1 vccd1 vccd1 _09878_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20350_ rbzero.debug_overlay.vplaneY\[-6\] rbzero.wall_tracer.rayAddendY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__xnor2_1
XFILLER_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19009_ _02665_ vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20281_ _03256_ vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__clkinv_2
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20617_ net84 _00633_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11350_ _03295_ _04051_ _04068_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__o21a_1
X_20548_ net123 _00564_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10301_ rbzero.tex_b1\[9\] rbzero.tex_b1\[10\] _03355_ vssd1 vssd1 vccd1 vccd1 _03360_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11281_ _03903_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__buf_4
XFILLER_197_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20479_ net94 _00495_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13020_ _05705_ _05708_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10232_ rbzero.tex_b1\[42\] rbzero.tex_b1\[43\] _03322_ vssd1 vssd1 vccd1 vccd1 _03324_
+ sky130_fd_sc_hd__mux2_1
XFILLER_234_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14971_ _07577_ _07583_ vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__nand2_1
XTAP_6799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16710_ rbzero.traced_texa\[10\] _09266_ _09267_ rbzero.wall_tracer.visualWallDist\[10\]
+ vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__a22o_1
X_13922_ _05651_ _06320_ _06472_ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__a21bo_1
XFILLER_43_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17690_ _09182_ _09978_ _01472_ _01473_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16641_ _09243_ vssd1 vssd1 vccd1 vccd1 _09247_ sky130_fd_sc_hd__clkbuf_4
XFILLER_235_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13853_ _06541_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__buf_2
XFILLER_169_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12804_ _05490_ _05492_ _05453_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__mux2_1
X_19360_ _02855_ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__buf_4
X_16572_ _09179_ _09180_ vssd1 vssd1 vccd1 vccd1 _09181_ sky130_fd_sc_hd__nor2_1
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13784_ _05662_ _06471_ _06472_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__a21boi_1
X_10996_ _03726_ vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__clkbuf_1
XFILLER_245_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18311_ rbzero.wall_tracer.trackDistY\[0\] rbzero.wall_tracer.stepDistY\[0\] _02072_
+ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__a21o_1
X_15523_ _07420_ _07421_ _07422_ _07645_ vssd1 vssd1 vccd1 vccd1 _08137_ sky130_fd_sc_hd__a211o_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12735_ _05361_ _05351_ _05422_ _05423_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__or4_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19291_ _02830_ vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18242_ _02015_ _02016_ _02017_ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__nand3_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _08067_ _08060_ vssd1 vssd1 vccd1 vccd1 _08068_ sky130_fd_sc_hd__or2_1
X_12666_ _05351_ _05354_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__nor2_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14405_ _06990_ _07064_ _07065_ vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__and3_1
X_11617_ _03910_ _04331_ _04332_ _04333_ _03945_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__o221a_1
XFILLER_204_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18173_ _01947_ _01952_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15385_ _07982_ _07998_ vssd1 vssd1 vccd1 vccd1 _07999_ sky130_fd_sc_hd__or2b_1
X_12597_ _05188_ _05285_ _03790_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__a21oi_1
XFILLER_141_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17124_ _08599_ _08510_ _08851_ _08979_ vssd1 vssd1 vccd1 vccd1 _09664_ sky130_fd_sc_hd__or4_1
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14336_ _05515_ _07024_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__nor2_1
X_11548_ rbzero.debug_overlay.vplaneY\[10\] _04236_ _04263_ _04265_ vssd1 vssd1 vccd1
+ vccd1 _04266_ sky130_fd_sc_hd__a211o_1
XFILLER_116_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17055_ _09592_ _09594_ _09595_ vssd1 vssd1 vccd1 vccd1 _09596_ sky130_fd_sc_hd__nand3_1
X_14267_ _06906_ _06954_ _06955_ _06903_ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__a211o_1
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11479_ _03802_ _03824_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__nand2_1
XFILLER_125_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16006_ _07672_ _07673_ _07400_ vssd1 vssd1 vccd1 vccd1 _08619_ sky130_fd_sc_hd__a21o_1
X_13218_ _05892_ _05899_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__xor2_1
XFILLER_174_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14198_ _06865_ _06866_ vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__xor2_1
XFILLER_174_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _05834_ _05836_ _05837_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__o21ai_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _01737_ _01738_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__xnor2_1
XFILLER_113_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16908_ _08478_ _08928_ vssd1 vssd1 vccd1 vccd1 _09450_ sky130_fd_sc_hd__and2_1
XFILLER_152_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17888_ _07619_ _07827_ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__nor2_1
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19627_ _02833_ _02995_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__nor2_1
X_16839_ _09379_ _09380_ vssd1 vssd1 vccd1 vccd1 _09381_ sky130_fd_sc_hd__nor2_1
XFILLER_96_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19558_ rbzero.pov.mosi rbzero.pov.mosi_buffer\[0\] _09243_ vssd1 vssd1 vccd1 vccd1
+ _02948_ sky130_fd_sc_hd__mux2_1
XFILLER_20_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18509_ _02238_ _02254_ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__xnor2_1
XFILLER_222_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19489_ _02912_ vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20402_ net121 _00433_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21382_ net113 _01398_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20333_ rbzero.debug_overlay.vplaneX\[-9\] rbzero.wall_tracer.rayAddendX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__or2_1
XFILLER_179_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20264_ _03255_ vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__clkinv_2
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20195_ rbzero.traced_texa\[4\] rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1 _03217_
+ sky130_fd_sc_hd__nor2_1
XFILLER_88_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10850_ _03650_ vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10781_ rbzero.tex_g0\[40\] rbzero.tex_g0\[39\] _03605_ vssd1 vssd1 vccd1 vccd1 _03614_
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12520_ _05162_ _05208_ _05161_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__o21ba_1
XFILLER_80_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ rbzero.debug_overlay.playerY\[4\] _05140_ _03798_ vssd1 vssd1 vccd1 vccd1
+ _05141_ sky130_fd_sc_hd__mux2_1
XFILLER_240_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11402_ rbzero.tex_r1\[49\] rbzero.tex_r1\[48\] _04119_ vssd1 vssd1 vccd1 vccd1 _04120_
+ sky130_fd_sc_hd__mux2_1
X_15170_ _07532_ _07585_ _07584_ vssd1 vssd1 vccd1 vccd1 _07784_ sky130_fd_sc_hd__a21o_1
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12382_ _05045_ _05074_ _05049_ _05034_ _05033_ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__a311o_2
XFILLER_240_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14121_ _06635_ _06808_ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__and2_1
X_11333_ rbzero.row_render.size\[7\] rbzero.row_render.size\[6\] vssd1 vssd1 vccd1
+ vccd1 _04052_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14052_ _06738_ _06739_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__xnor2_1
XFILLER_180_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11264_ _03924_ _03977_ _03982_ _03899_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__a211o_1
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13003_ _05565_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__buf_2
X_10215_ rbzero.tex_b1\[50\] rbzero.tex_b1\[51\] _03311_ vssd1 vssd1 vccd1 vccd1 _03315_
+ sky130_fd_sc_hd__mux2_1
XFILLER_234_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18860_ rbzero.spi_registers.sclk_buffer\[2\] rbzero.spi_registers.sclk_buffer\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__and2b_1
XTAP_6530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11195_ _03860_ _03894_ _03907_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__or3b_2
XTAP_6541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17811_ _01593_ _01594_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__and2b_1
XTAP_6552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18791_ _02508_ _02511_ _02507_ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__a21o_1
XTAP_6585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17742_ _01469_ _01450_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__and2b_1
XTAP_5873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14954_ _07213_ _07164_ _07346_ vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__a21o_1
XFILLER_153_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13905_ _06310_ _06389_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__nor2_1
X_17673_ _08923_ _09470_ _08240_ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__a21o_1
X_14885_ _03794_ _05114_ _07498_ vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__or3_1
XFILLER_223_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19412_ rbzero.pov.spi_buffer\[4\] rbzero.pov.spi_buffer\[5\] _02866_ vssd1 vssd1
+ vccd1 vccd1 _02872_ sky130_fd_sc_hd__mux2_1
X_16624_ _09231_ _09229_ vssd1 vssd1 vccd1 vccd1 _09233_ sky130_fd_sc_hd__or2b_1
X_13836_ _06465_ _06523_ _06522_ vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__a21o_1
XFILLER_1_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19343_ _02857_ vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__clkinv_2
XFILLER_90_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16555_ _07805_ _07685_ _07712_ _08067_ vssd1 vssd1 vccd1 vccd1 _09164_ sky130_fd_sc_hd__o22a_1
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13767_ _06430_ _06448_ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__xnor2_1
X_10979_ rbzero.tex_b0\[10\] rbzero.tex_b0\[9\] _03715_ vssd1 vssd1 vccd1 vccd1 _03718_
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15506_ _08118_ _08119_ vssd1 vssd1 vccd1 vccd1 _08120_ sky130_fd_sc_hd__nor2_1
XFILLER_206_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12718_ _05405_ _05406_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__or2b_1
X_19274_ _02821_ vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__clkbuf_1
X_16486_ _08955_ _09095_ vssd1 vssd1 vccd1 vccd1 _09096_ sky130_fd_sc_hd__xor2_4
X_13698_ _06165_ _06175_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__nand2_1
XFILLER_143_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18225_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.stepDistY\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__or2_1
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15437_ _08042_ _08044_ vssd1 vssd1 vccd1 vccd1 _08051_ sky130_fd_sc_hd__xor2_1
XFILLER_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12649_ _05336_ _05337_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__nor2_1
XFILLER_54_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18156_ _01882_ _01884_ _01935_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__o21a_1
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15368_ _07980_ _07963_ vssd1 vssd1 vccd1 vccd1 _07982_ sky130_fd_sc_hd__xor2_1
XFILLER_172_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17107_ _09303_ _09645_ _09647_ _09282_ vssd1 vssd1 vccd1 vccd1 _09648_ sky130_fd_sc_hd__a31o_1
X_14319_ _06962_ _06964_ vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__and2_1
XFILLER_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18087_ _01865_ _01867_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__nor2_1
XFILLER_171_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15299_ _07911_ _07912_ vssd1 vssd1 vccd1 vccd1 _07913_ sky130_fd_sc_hd__nor2_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17038_ _07805_ _07834_ vssd1 vssd1 vccd1 vccd1 _09579_ sky130_fd_sc_hd__or2_1
XFILLER_172_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ rbzero.pov.spi_buffer\[42\] rbzero.pov.ready_buffer\[42\] _02651_ vssd1 vssd1
+ vccd1 vccd1 _02655_ sky130_fd_sc_hd__mux2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20951_ net76 _00967_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_54_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20882_ net58 _00898_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21365_ _00388_ _01381_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20316_ rbzero.traced_texVinit\[6\] _09266_ _09099_ _09261_ vssd1 vssd1 vccd1 vccd1
+ _01400_ sky130_fd_sc_hd__a22o_1
XFILLER_135_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21296_ net134 _01312_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20247_ _03253_ vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__clkinv_2
XFILLER_192_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20178_ _03202_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__inv_2
XFILLER_49_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11951_ _04650_ _04651_ _04661_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__a21o_1
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10902_ _03677_ vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__clkbuf_1
X_14670_ rbzero.wall_tracer.stepDistX\[-10\] _07147_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _07309_ sky130_fd_sc_hd__mux2_1
XFILLER_166_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11882_ rbzero.row_render.wall\[0\] vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__inv_2
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13621_ _05746_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__buf_2
X_10833_ _03641_ vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16340_ _08746_ _08813_ _08950_ vssd1 vssd1 vccd1 vccd1 _08951_ sky130_fd_sc_hd__a21oi_1
XFILLER_186_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13552_ _06239_ _06240_ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__and2_1
XFILLER_164_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10764_ _03604_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__clkbuf_4
XFILLER_207_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12503_ _05188_ _05191_ _03790_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__a21o_1
XFILLER_125_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16271_ _08759_ _08761_ vssd1 vssd1 vccd1 vccd1 _08882_ sky130_fd_sc_hd__nor2_1
XFILLER_186_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13483_ _06171_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__buf_2
XFILLER_16_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10695_ rbzero.tex_g1\[16\] rbzero.tex_g1\[17\] _03563_ vssd1 vssd1 vccd1 vccd1 _03569_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18010_ _01789_ _01791_ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__nor2_1
XFILLER_51_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15222_ _07834_ _07835_ _07663_ _07680_ vssd1 vssd1 vccd1 vccd1 _07836_ sky130_fd_sc_hd__or4_1
XFILLER_185_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12434_ _05124_ _05125_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__or2_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15153_ _04929_ _07698_ _07651_ _07765_ vssd1 vssd1 vccd1 vccd1 _07767_ sky130_fd_sc_hd__a31o_1
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12365_ rbzero.debug_overlay.facingY\[-1\] rbzero.wall_tracer.rayAddendY\[7\] _05057_
+ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__a21oi_1
XFILLER_181_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14104_ _06791_ _06792_ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__nor2_1
X_11316_ rbzero.floor_leak\[2\] _03945_ _03949_ rbzero.floor_leak\[3\] _04034_ vssd1
+ vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__o221a_1
XFILLER_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15084_ rbzero.wall_tracer.visualWallDist\[-12\] _03794_ vssd1 vssd1 vccd1 vccd1
+ _07698_ sky130_fd_sc_hd__and2_4
X_19961_ _03119_ vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__clkinv_2
X_12296_ _04982_ _04988_ _04989_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__or3_1
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14035_ _06717_ _06718_ _06722_ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__nand3_1
X_18912_ _02614_ vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__clkbuf_1
XTAP_7050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11247_ rbzero.tex_r0\[47\] _03964_ _03965_ _03930_ vssd1 vssd1 vccd1 vccd1 _03966_
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19892_ _02862_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__buf_4
XTAP_7061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18843_ _02428_ rbzero.debug_overlay.vplaneY\[-1\] _02552_ _02510_ vssd1 vssd1 vccd1
+ vccd1 _02561_ sky130_fd_sc_hd__a211oi_1
XTAP_6360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11178_ _03867_ _03846_ _03864_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__nor3_1
XFILLER_132_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18774_ _02495_ _02496_ _03812_ vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__o21ai_1
XFILLER_212_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15986_ _08296_ vssd1 vssd1 vccd1 vccd1 _08599_ sky130_fd_sc_hd__buf_2
XTAP_5670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17725_ _01507_ _01508_ _01509_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__or3_1
XTAP_5692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14937_ _07423_ _07485_ _07542_ _07550_ vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__or4_1
XFILLER_36_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17656_ _01438_ _01440_ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__nor2_1
X_14868_ _07349_ rbzero.wall_tracer.stepDistY\[-7\] rbzero.wall_tracer.state\[6\]
+ vssd1 vssd1 vccd1 vccd1 _07482_ sky130_fd_sc_hd__a21oi_2
XFILLER_169_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16607_ _09214_ _09215_ vssd1 vssd1 vccd1 vccd1 _09216_ sky130_fd_sc_hd__xor2_1
XFILLER_224_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13819_ _06476_ _06475_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__and2_1
XFILLER_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17587_ _09989_ _09990_ _09991_ vssd1 vssd1 vccd1 vccd1 _10124_ sky130_fd_sc_hd__nand3_1
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14799_ _07411_ _07412_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__nand2_1
XFILLER_95_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19326_ _04702_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__buf_4
X_16538_ _09143_ _09146_ vssd1 vssd1 vccd1 vccd1 _09147_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19257_ rbzero.spi_registers.spi_done _03292_ _02582_ vssd1 vssd1 vccd1 vccd1 _02812_
+ sky130_fd_sc_hd__and3_1
X_16469_ _08941_ _08943_ vssd1 vssd1 vccd1 vccd1 _09079_ sky130_fd_sc_hd__nand2_1
X_18208_ _01911_ _01915_ _01987_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__o21a_1
XFILLER_176_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19188_ rbzero.spi_registers.new_floor\[5\] rbzero.spi_registers.got_new_floor _02724_
+ _02753_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__a31o_1
XFILLER_191_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18139_ _01825_ _01918_ _01917_ _09351_ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__a31o_1
XFILLER_145_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21150_ _00199_ _01166_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20101_ rbzero.traced_texa\[-11\] rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1 _03138_
+ sky130_fd_sc_hd__or2_1
XFILLER_160_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21081_ _00130_ _01097_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20032_ _03126_ vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__clkinv_2
XFILLER_140_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20934_ net69 _00950_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[71\] sky130_fd_sc_hd__dfxtp_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20865_ net79 _00881_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20796_ net84 _00812_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_210_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10480_ rbzero.tex_r0\[55\] rbzero.tex_r0\[54\] _03446_ vssd1 vssd1 vccd1 vccd1 _03456_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12150_ _04830_ _04855_ _04856_ _04844_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__a22o_1
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21348_ _00371_ _01364_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11101_ gpout0.vpos\[9\] gpout0.vpos\[8\] gpout0.vpos\[7\] net2 vssd1 vssd1 vccd1
+ vccd1 _03820_ sky130_fd_sc_hd__or4b_1
XFILLER_11_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12081_ _04773_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__inv_2
XFILLER_150_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21279_ _00328_ _01295_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11032_ rbzero.map_rom.f4 _03733_ _03758_ _03759_ vssd1 vssd1 vccd1 vccd1 _03760_
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15840_ _08450_ _08452_ _08453_ vssd1 vssd1 vccd1 vccd1 _08454_ sky130_fd_sc_hd__a21o_1
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15771_ _08382_ _08384_ vssd1 vssd1 vccd1 vccd1 _08385_ sky130_fd_sc_hd__nor2_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12983_ _05447_ _05479_ _05482_ _05487_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__o22ai_4
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17510_ _09906_ _10046_ vssd1 vssd1 vccd1 vccd1 _10047_ sky130_fd_sc_hd__xnor2_1
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14722_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__buf_4
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18490_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.debug_overlay.vplaneX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__and2_1
X_11934_ net48 _04611_ _04618_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__and3_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _09449_ _09978_ _09851_ vssd1 vssd1 vccd1 vccd1 _09979_ sky130_fd_sc_hd__or3_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14653_ rbzero.wall_tracer.visualWallDist\[7\] _07252_ vssd1 vssd1 vccd1 vccd1 _07299_
+ sky130_fd_sc_hd__or2_1
XFILLER_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ rbzero.tex_b1\[7\] rbzero.tex_b1\[6\] _04544_ vssd1 vssd1 vccd1 vccd1 _04579_
+ sky130_fd_sc_hd__mux2_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _05434_ _05847_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__or2_1
XFILLER_60_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17372_ _09901_ _09902_ _09908_ vssd1 vssd1 vccd1 vccd1 _09910_ sky130_fd_sc_hd__and3_1
X_10816_ _03632_ vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__clkbuf_1
X_14584_ _07248_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__clkbuf_4
X_11796_ rbzero.tex_b0\[10\] _03936_ _03929_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__a21o_1
XFILLER_92_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19111_ _02722_ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__buf_2
X_16323_ _08794_ _08795_ vssd1 vssd1 vccd1 vccd1 _08934_ sky130_fd_sc_hd__and2b_1
X_13535_ _06218_ _06220_ _06223_ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__a21o_1
XFILLER_159_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10747_ rbzero.tex_g0\[56\] rbzero.tex_g0\[55\] _03593_ vssd1 vssd1 vccd1 vccd1 _03596_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19042_ _02682_ vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16254_ _08592_ _08296_ _07621_ rbzero.wall_tracer.visualWallDist\[4\] vssd1 vssd1
+ vccd1 vccd1 _08865_ sky130_fd_sc_hd__or4b_1
X_13466_ _06148_ _06150_ _06153_ _06154_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__a31o_1
XFILLER_139_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10678_ rbzero.tex_g1\[24\] rbzero.tex_g1\[25\] _03552_ vssd1 vssd1 vccd1 vccd1 _03560_
+ sky130_fd_sc_hd__mux2_1
XFILLER_220_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15205_ _07101_ _07220_ vssd1 vssd1 vccd1 vccd1 _07819_ sky130_fd_sc_hd__and2_1
X_12417_ _05108_ _05109_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__nor2_1
X_16185_ _07847_ _08634_ vssd1 vssd1 vccd1 vccd1 _08797_ sky130_fd_sc_hd__nor2_1
XFILLER_182_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13397_ _06070_ _06082_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__xor2_1
XFILLER_160_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15136_ _07748_ _07743_ _07749_ vssd1 vssd1 vccd1 vccd1 _07750_ sky130_fd_sc_hd__o21ai_1
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12348_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] _05039_
+ _05040_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__a31o_1
XFILLER_245_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15067_ _07472_ _07680_ _07674_ vssd1 vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__or3_1
X_12279_ _04967_ _04971_ _04972_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__a21o_1
X_19944_ _03117_ vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__clkinv_2
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14018_ _06658_ _06678_ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19875_ _03110_ vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__clkinv_2
XFILLER_68_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18826_ _02528_ _02533_ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__nand2_1
XFILLER_110_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18757_ _02479_ _02480_ vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__nor2_1
XFILLER_243_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15969_ _08567_ _08582_ vssd1 vssd1 vccd1 vccd1 _08583_ sky130_fd_sc_hd__xor2_1
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17708_ _01491_ _01492_ vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__and2b_1
XFILLER_224_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18688_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__or2_1
XFILLER_247_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17639_ _10173_ _10174_ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__or2_1
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20650_ net63 _00666_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_210_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19309_ _02837_ _02843_ _02838_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__a21boi_1
XFILLER_210_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20581_ net93 _00597_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21202_ _00251_ _01218_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21133_ _00182_ _01149_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21064_ _00113_ _01080_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20015_ _03124_ vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__clkinv_2
XFILLER_189_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20917_ net68 _00933_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[54\] sky130_fd_sc_hd__dfxtp_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11650_ _03910_ _04364_ _04365_ _04366_ _03945_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__o221a_1
XFILLER_202_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20848_ _00066_ _00864_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10601_ rbzero.tex_g1\[61\] rbzero.tex_g1\[62\] _03519_ vssd1 vssd1 vccd1 vccd1 _03520_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout63 net64 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11581_ _04276_ _04298_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__nand2_1
Xfanout74 net77 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__buf_2
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20779_ net88 _00795_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout85 net86 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13320_ _05625_ _06008_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__nand2_1
Xfanout96 net97 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__buf_2
X_10532_ _03483_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13251_ _05615_ _05939_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10463_ _03447_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12202_ net42 _04885_ _04907_ net36 vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13182_ _05856_ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10394_ rbzero.tex_r1\[29\] rbzero.tex_r1\[30\] _03400_ vssd1 vssd1 vccd1 vccd1 _03409_
+ sky130_fd_sc_hd__mux2_1
X_12133_ _04825_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__inv_2
XFILLER_237_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17990_ _01770_ _01771_ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16941_ _09206_ _09213_ _09482_ vssd1 vssd1 vccd1 vccd1 _09483_ sky130_fd_sc_hd__a21o_1
X_12064_ _04768_ o_rgb[7] _04771_ net25 vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__a211o_1
XFILLER_78_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11015_ rbzero.map_rom.d6 vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__inv_2
X_19660_ rbzero.pov.ready_buffer\[49\] _02958_ _03008_ _03023_ vssd1 vssd1 vccd1 vccd1
+ _03024_ sky130_fd_sc_hd__a211o_1
X_16872_ _09017_ _09021_ _09147_ vssd1 vssd1 vccd1 vccd1 _09414_ sky130_fd_sc_hd__a21oi_1
XFILLER_133_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18611_ rbzero.map_rom.f3 _07491_ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15823_ _08409_ _08404_ vssd1 vssd1 vccd1 vccd1 _08437_ sky130_fd_sc_hd__or2_1
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19591_ _07394_ _02960_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__nand2_1
XFILLER_133_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ _03819_ _02284_ _02285_ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__nor3_1
X_15754_ _07529_ _07984_ _07646_ vssd1 vssd1 vccd1 vccd1 _08368_ sky130_fd_sc_hd__a21o_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12966_ _05621_ _05638_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__nor2_1
XFILLER_161_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14705_ rbzero.wall_tracer.stepDistX\[7\] _07229_ _04931_ vssd1 vssd1 vccd1 vccd1
+ _07327_ sky130_fd_sc_hd__mux2_1
XFILLER_166_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ gpout0.vpos\[2\] vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__buf_2
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18473_ _02204_ _02218_ _02219_ _02220_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__nand4_2
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15685_ _08294_ _08297_ _08298_ vssd1 vssd1 vccd1 vccd1 _08299_ sky130_fd_sc_hd__a21bo_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _05462_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__clkbuf_4
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17424_ _08240_ _09055_ vssd1 vssd1 vccd1 vccd1 _09962_ sky130_fd_sc_hd__or2b_1
XFILLER_178_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ rbzero.wall_tracer.visualWallDist\[2\] _07252_ vssd1 vssd1 vccd1 vccd1 _07287_
+ sky130_fd_sc_hd__or2_1
XFILLER_127_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11848_ rbzero.tex_b1\[25\] rbzero.tex_b1\[24\] _03934_ vssd1 vssd1 vccd1 vccd1 _04562_
+ sky130_fd_sc_hd__mux2_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17355_ _09303_ _09892_ _09893_ _09282_ vssd1 vssd1 vccd1 vccd1 _09894_ sky130_fd_sc_hd__a31o_1
X_14567_ _07235_ vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11779_ rbzero.tex_b0\[22\] _03962_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__and2_1
XFILLER_201_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16306_ _08916_ vssd1 vssd1 vccd1 vccd1 _08917_ sky130_fd_sc_hd__clkbuf_4
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13518_ _06195_ _06206_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__xnor2_1
X_17286_ _09789_ _09824_ vssd1 vssd1 vccd1 vccd1 _09825_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14498_ rbzero.wall_tracer.stepDistY\[-6\] _07180_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _07181_ sky130_fd_sc_hd__mux2_1
XFILLER_105_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19025_ rbzero.pov.spi_buffer\[59\] rbzero.pov.ready_buffer\[59\] _02673_ vssd1 vssd1
+ vccd1 vccd1 _02674_ sky130_fd_sc_hd__mux2_1
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16237_ _08766_ _08747_ vssd1 vssd1 vccd1 vccd1 _08848_ sky130_fd_sc_hd__or2b_1
X_13449_ _06133_ _06131_ _06137_ _06122_ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__a211o_1
XFILLER_127_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16168_ _07696_ _08640_ vssd1 vssd1 vccd1 vccd1 _08780_ sky130_fd_sc_hd__and2_2
XFILLER_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15119_ _07730_ _07732_ _07351_ vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__a21oi_1
XFILLER_114_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16099_ _08693_ _08695_ vssd1 vssd1 vccd1 vccd1 _08711_ sky130_fd_sc_hd__nor2_1
XFILLER_47_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19927_ _03116_ vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__clkinv_2
XFILLER_151_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19858_ _03108_ vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__clkinv_2
XFILLER_64_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18809_ _02509_ rbzero.wall_tracer.rayAddendY\[7\] vssd1 vssd1 vccd1 vccd1 _02529_
+ sky130_fd_sc_hd__or2_1
XFILLER_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19789_ _09245_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__clkbuf_4
XFILLER_110_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20702_ net87 _00718_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20633_ net54 _00649_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20564_ net123 _00580_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20495_ net127 _00511_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21116_ _00165_ _01132_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_6937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21047_ _00096_ _01063_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12820_ _05508_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__inv_2
XFILLER_74_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _05361_ _05363_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__nor2_2
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ rbzero.tex_g1\[49\] rbzero.tex_g1\[48\] _04378_ vssd1 vssd1 vccd1 vccd1 _04418_
+ sky130_fd_sc_hd__mux2_1
XFILLER_231_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15470_ _08082_ _08083_ vssd1 vssd1 vccd1 vccd1 _08084_ sky130_fd_sc_hd__xor2_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12682_ _05261_ _05249_ _05295_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__o21a_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14421_ _05527_ _07106_ _07109_ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__a21oi_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _03957_ _04347_ _04348_ _04349_ _03945_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__o221a_1
XFILLER_230_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17140_ _07619_ _07709_ vssd1 vssd1 vccd1 vccd1 _09680_ sky130_fd_sc_hd__nor2_1
X_14352_ _07039_ _07040_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__or2b_1
XFILLER_156_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11564_ _04229_ _04201_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__nor2_1
XFILLER_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13303_ _05983_ _05989_ _05991_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__o21a_1
X_17071_ _09476_ _09608_ _09609_ _09611_ vssd1 vssd1 vccd1 vccd1 _09612_ sky130_fd_sc_hd__and4b_1
X_10515_ _03474_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__clkbuf_1
X_14283_ _06629_ _06971_ _06573_ vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__a21oi_1
XFILLER_196_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11495_ _04203_ _04212_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__nor2_1
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16022_ _07826_ _07471_ _08628_ _08634_ vssd1 vssd1 vccd1 vccd1 _08635_ sky130_fd_sc_hd__or4_1
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13234_ _05921_ _05909_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__and2b_1
X_10446_ _03436_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13165_ _05846_ _05853_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10377_ _03388_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__clkbuf_4
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12116_ _04820_ _04118_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__nor2_1
X_17973_ _01625_ _01645_ _01623_ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__a21oi_2
X_13096_ _05682_ _05683_ _05684_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__a21oi_1
XFILLER_124_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16924_ _08398_ _09200_ _07826_ vssd1 vssd1 vccd1 vccd1 _09466_ sky130_fd_sc_hd__o21ai_1
X_12047_ net52 _04717_ _04718_ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__and3_1
X_19712_ rbzero.pov.ready_buffer\[34\] _03061_ _03063_ rbzero.debug_overlay.facingX\[-8\]
+ _03064_ vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__a221o_1
XFILLER_242_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16855_ _08510_ _08985_ _09130_ _09131_ vssd1 vssd1 vccd1 vccd1 _09397_ sky130_fd_sc_hd__o31a_1
X_19643_ _03008_ _03010_ _03011_ _02978_ vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__o211a_1
XFILLER_66_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15806_ _07835_ _08059_ _08393_ vssd1 vssd1 vccd1 vccd1 _08420_ sky130_fd_sc_hd__o21bai_1
XFILLER_4_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19574_ _02834_ vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__buf_2
X_16786_ rbzero.wall_tracer.trackDistX\[-5\] rbzero.wall_tracer.stepDistX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _09333_ sky130_fd_sc_hd__nand2_1
XFILLER_225_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13998_ _06575_ _06627_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__and2_1
XFILLER_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18525_ _09256_ _02269_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__nand2_1
X_15737_ _08323_ _08350_ vssd1 vssd1 vccd1 vccd1 _08351_ sky130_fd_sc_hd__or2_1
XFILLER_98_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12949_ _05637_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__buf_2
XFILLER_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18456_ rbzero.debug_overlay.vplaneX\[0\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__nand2_1
X_15668_ _08272_ _08060_ _08234_ _08280_ _08281_ vssd1 vssd1 vccd1 vccd1 _08282_ sky130_fd_sc_hd__o41a_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17407_ _09932_ _09943_ vssd1 vssd1 vccd1 vccd1 _09945_ sky130_fd_sc_hd__or2_1
X_14619_ rbzero.wall_tracer.trackDistY\[-3\] vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__inv_2
XFILLER_18_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18387_ rbzero.spi_registers.new_vinf rbzero.spi_registers.spi_buffer\[0\] _02141_
+ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__mux2_1
X_15599_ _08192_ _08211_ vssd1 vssd1 vccd1 vccd1 _08213_ sky130_fd_sc_hd__or2b_1
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17338_ _09874_ _09876_ vssd1 vssd1 vccd1 vccd1 _09877_ sky130_fd_sc_hd__xor2_1
XFILLER_18_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17269_ _09681_ _09685_ _09682_ vssd1 vssd1 vccd1 vccd1 _09808_ sky130_fd_sc_hd__a21bo_1
XFILLER_146_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19008_ rbzero.pov.spi_buffer\[51\] rbzero.pov.ready_buffer\[51\] _02662_ vssd1 vssd1
+ vccd1 vccd1 _02665_ sky130_fd_sc_hd__mux2_1
XFILLER_106_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20280_ _03256_ vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__clkinv_2
XFILLER_179_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20616_ net99 _00632_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20547_ net125 _00563_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10300_ _03359_ vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11280_ rbzero.tex_r0\[29\] rbzero.tex_r0\[28\] _03936_ vssd1 vssd1 vccd1 vccd1 _03999_
+ sky130_fd_sc_hd__mux2_1
X_20478_ net94 _00494_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10231_ _03323_ vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_238_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14970_ _07577_ _07583_ vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__nor2_1
XTAP_6789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13921_ _06516_ _06517_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__xnor2_1
XFILLER_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16640_ _09246_ vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__clkbuf_1
X_13852_ _06173_ _06540_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__nand2_1
XFILLER_210_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ _05491_ _05423_ _05429_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__mux2_1
X_16571_ _09161_ _09178_ vssd1 vssd1 vccd1 vccd1 _09180_ sky130_fd_sc_hd__nor2_1
XFILLER_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13783_ _06260_ _06289_ _06303_ _06470_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__a211o_1
XFILLER_204_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10995_ rbzero.tex_b0\[2\] rbzero.tex_b0\[1\] _03445_ vssd1 vssd1 vccd1 vccd1 _03726_
+ sky130_fd_sc_hd__mux2_1
X_18310_ rbzero.wall_tracer.trackDistY\[1\] rbzero.wall_tracer.stepDistY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__nand2_1
XFILLER_43_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15522_ _07466_ _07664_ vssd1 vssd1 vccd1 vccd1 _08136_ sky130_fd_sc_hd__nor2_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ _05333_ _05334_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__nor2_1
X_19290_ rbzero.spi_registers.new_vshift\[4\] rbzero.spi_registers.spi_buffer\[4\]
+ _02825_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__mux2_1
XFILLER_245_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18241_ _02008_ _02009_ _02010_ vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__o21bai_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _07591_ vssd1 vssd1 vccd1 vccd1 _08067_ sky130_fd_sc_hd__clkbuf_4
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12665_ _05353_ _05335_ _05343_ _05346_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__or4_1
XFILLER_54_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14404_ _06990_ _06986_ _06989_ vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__and3_1
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18172_ _01950_ _01951_ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__xor2_1
XFILLER_180_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11616_ rbzero.tex_g0\[10\] _03974_ _03929_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__a21o_1
XFILLER_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15384_ _07610_ _07983_ _07990_ _07997_ vssd1 vssd1 vccd1 vccd1 _07998_ sky130_fd_sc_hd__o31ai_1
XFILLER_50_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12596_ rbzero.wall_tracer.visualWallDist\[6\] _05190_ vssd1 vssd1 vccd1 vccd1 _05285_
+ sky130_fd_sc_hd__nand2_1
X_17123_ _08599_ _08852_ _09373_ _08510_ vssd1 vssd1 vccd1 vccd1 _09663_ sky130_fd_sc_hd__o22ai_1
XFILLER_204_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14335_ _06959_ _06961_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__xnor2_4
XFILLER_15_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11547_ rbzero.debug_overlay.vplaneY\[-9\] _04240_ _04218_ rbzero.debug_overlay.vplaneY\[-8\]
+ _04264_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__a221o_1
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17054_ _07858_ _08917_ vssd1 vssd1 vccd1 vccd1 _09595_ sky130_fd_sc_hd__nor2_1
XFILLER_167_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14266_ _06885_ _06905_ vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__nor2_1
XFILLER_183_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11478_ _03806_ _04195_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__or2_1
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16005_ _07472_ _07641_ _07379_ vssd1 vssd1 vccd1 vccd1 _08618_ sky130_fd_sc_hd__a21o_1
X_13217_ _05802_ _05813_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__xnor2_1
X_10429_ _03427_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__clkbuf_1
X_14197_ _06855_ _06872_ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13148_ _05832_ _05833_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__nand2_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17956_ _09428_ _08787_ vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__nor2_1
X_13079_ _05607_ _05767_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__nor2_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16907_ _07400_ vssd1 vssd1 vccd1 vccd1 _09449_ sky130_fd_sc_hd__buf_2
X_17887_ _01568_ _01571_ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__nand2_1
XFILLER_22_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19626_ rbzero.debug_overlay.playerX\[3\] _02960_ _02997_ _02989_ vssd1 vssd1 vccd1
+ vccd1 _00972_ sky130_fd_sc_hd__a211o_1
X_16838_ _09156_ _09372_ _09378_ vssd1 vssd1 vccd1 vccd1 _09380_ sky130_fd_sc_hd__and3_1
XFILLER_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16769_ rbzero.wall_tracer.trackDistX\[-7\] rbzero.wall_tracer.stepDistX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _09318_ sky130_fd_sc_hd__or2_1
X_19557_ _02947_ vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__clkbuf_1
XFILLER_241_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18508_ _02252_ _02253_ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__xnor2_1
X_19488_ rbzero.pov.spi_buffer\[40\] rbzero.pov.spi_buffer\[41\] _02910_ vssd1 vssd1
+ vccd1 vccd1 _02912_ sky130_fd_sc_hd__mux2_1
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18439_ rbzero.wall_tracer.rayAddendX\[-2\] _00013_ _02186_ _02189_ vssd1 vssd1 vccd1
+ vccd1 _00593_ sky130_fd_sc_hd__o22a_1
XFILLER_210_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20401_ net121 _00432_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-10\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_33_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21381_ net97 _01397_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20332_ _03266_ vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20263_ _03255_ vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__clkinv_2
XFILLER_89_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20194_ _03211_ _03213_ _03212_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__a21boi_1
XFILLER_192_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _03613_ vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12450_ _05138_ _05139_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__xnor2_1
XFILLER_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11401_ _03934_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__clkbuf_4
XFILLER_166_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12381_ _05044_ _05043_ _05047_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__nand3_1
XFILLER_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14120_ _06635_ _06808_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__nor2_1
XFILLER_126_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11332_ rbzero.row_render.size\[9\] _04048_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__nor2_1
XFILLER_197_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14051_ _06738_ _06739_ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__nand2_1
XFILLER_181_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11263_ _03932_ _03978_ _03979_ _03981_ _03946_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__o221a_1
XFILLER_238_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13002_ _05688_ _05690_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10214_ _03314_ vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11194_ rbzero.tex_r0\[53\] rbzero.tex_r0\[52\] _03904_ vssd1 vssd1 vccd1 vccd1 _03913_
+ sky130_fd_sc_hd__mux2_1
XTAP_6520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17810_ _01590_ _01592_ vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__nand2_1
XTAP_6553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18790_ _02507_ _02508_ _02511_ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__nand3_1
XTAP_5830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17741_ _01429_ _01443_ _01441_ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__a21o_1
XTAP_5852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14953_ _07566_ vssd1 vssd1 vccd1 vccd1 _07567_ sky130_fd_sc_hd__buf_2
XTAP_5874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13904_ _06590_ _06592_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__xnor2_1
X_17672_ _01455_ _01456_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__and2_1
XFILLER_247_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14884_ rbzero.debug_overlay.playerY\[-1\] rbzero.debug_overlay.playerY\[-2\] _07497_
+ vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__or3_1
XFILLER_1_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16623_ _09229_ _09231_ vssd1 vssd1 vccd1 vccd1 _09232_ sky130_fd_sc_hd__and2b_1
X_19411_ _02871_ vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__clkbuf_1
X_13835_ _06465_ _06522_ _06523_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__nand3_1
XFILLER_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16554_ _07793_ vssd1 vssd1 vccd1 vccd1 _09163_ sky130_fd_sc_hd__buf_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19342_ _02857_ vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__clkinv_2
X_13766_ _06453_ _06454_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__and2_1
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10978_ _03717_ vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__clkbuf_1
X_15505_ _07399_ _07508_ _07575_ _07378_ vssd1 vssd1 vccd1 vccd1 _08119_ sky130_fd_sc_hd__o22a_1
XFILLER_241_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12717_ _05399_ _05404_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__nand2_2
X_19273_ rbzero.spi_registers.new_other\[8\] rbzero.spi_registers.spi_buffer\[8\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__mux2_1
XFILLER_231_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16485_ _08844_ _09094_ vssd1 vssd1 vccd1 vccd1 _09095_ sky130_fd_sc_hd__xor2_2
X_13697_ _05767_ _06331_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__or2_1
XFILLER_182_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18224_ rbzero.wall_tracer.trackDistY\[-12\] _01996_ _02002_ _09278_ vssd1 vssd1
+ vccd1 vccd1 _00565_ sky130_fd_sc_hd__o22a_1
XFILLER_248_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15436_ _08045_ _08047_ _08048_ _08049_ vssd1 vssd1 vccd1 vccd1 _08050_ sky130_fd_sc_hd__o22a_1
X_12648_ _05227_ _05229_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__and2_2
XFILLER_50_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18155_ _01871_ _01885_ vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__or2b_1
XFILLER_200_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15367_ _07963_ _07980_ vssd1 vssd1 vccd1 vccd1 _07981_ sky130_fd_sc_hd__or2b_1
XFILLER_117_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12579_ _05108_ _05109_ _03815_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__o21ai_1
XFILLER_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17106_ _09646_ vssd1 vssd1 vccd1 vccd1 _09647_ sky130_fd_sc_hd__inv_2
XFILLER_89_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14318_ _05569_ vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__clkbuf_2
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18086_ _09833_ _08725_ _01769_ _01866_ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__o31a_1
X_15298_ _07616_ _07617_ _07621_ _07788_ vssd1 vssd1 vccd1 vccd1 _07912_ sky130_fd_sc_hd__o22a_1
XFILLER_183_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17037_ _09170_ _09576_ _09577_ _09434_ vssd1 vssd1 vccd1 vccd1 _09578_ sky130_fd_sc_hd__o22ai_2
XFILLER_172_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14249_ _06799_ _06937_ vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__nand2_1
XFILLER_176_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18988_ _02654_ vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__clkbuf_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ rbzero.wall_tracer.trackDistX\[8\] rbzero.wall_tracer.stepDistX\[8\] vssd1
+ vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__nor2_1
XFILLER_26_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20950_ net76 _00966_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19609_ _02982_ _02983_ _02835_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__a21oi_1
XFILLER_148_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20881_ net55 _00897_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_226_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21364_ _00387_ _01380_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20315_ rbzero.traced_texVinit\[5\] _09266_ _08959_ _09261_ vssd1 vssd1 vccd1 vccd1
+ _01399_ sky130_fd_sc_hd__a22o_1
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21295_ net134 _01311_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20246_ _03253_ vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__clkinv_2
XFILLER_157_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20177_ _03199_ _03200_ _03201_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__and3_1
XFILLER_190_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ _04630_ net11 _04657_ _04660_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__a31o_1
XFILLER_229_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ rbzero.tex_b0\[47\] rbzero.tex_b0\[46\] _03671_ vssd1 vssd1 vccd1 vccd1 _03677_
+ sky130_fd_sc_hd__mux2_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11881_ _04592_ rbzero.row_render.wall\[1\] _03288_ vssd1 vssd1 vccd1 vccd1 _04594_
+ sky130_fd_sc_hd__o21a_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13620_ _06230_ _06306_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__nand2_1
XFILLER_246_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10832_ rbzero.tex_g0\[16\] rbzero.tex_g0\[15\] _03638_ vssd1 vssd1 vccd1 vccd1 _03641_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13551_ _05645_ _05624_ _05701_ _05692_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__a22o_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10763_ _03444_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__clkbuf_4
XFILLER_186_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12502_ rbzero.wall_tracer.visualWallDist\[9\] _05190_ vssd1 vssd1 vccd1 vccd1 _05191_
+ sky130_fd_sc_hd__nand2_1
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16270_ _08847_ _08880_ vssd1 vssd1 vccd1 vccd1 _08881_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13482_ _06169_ _06170_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__or2_1
XFILLER_157_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10694_ _03568_ vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15221_ _07646_ vssd1 vssd1 vccd1 vccd1 _07835_ sky130_fd_sc_hd__buf_4
X_12433_ rbzero.map_rom.d6 _05117_ _05115_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__a21o_1
XFILLER_240_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15152_ _04929_ _07698_ _07651_ _07765_ vssd1 vssd1 vccd1 vccd1 _07766_ sky130_fd_sc_hd__and4_1
XFILLER_51_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12364_ rbzero.debug_overlay.facingY\[0\] rbzero.wall_tracer.rayAddendY\[8\] vssd1
+ vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__and2_1
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14103_ _06786_ _06790_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__nor2_1
XFILLER_5_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11315_ rbzero.floor_leak\[1\] _03928_ _03944_ rbzero.floor_leak\[2\] _04033_ vssd1
+ vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__a221o_1
X_15083_ _07434_ vssd1 vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__clkinv_4
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19960_ _03119_ vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__clkinv_2
X_12295_ _04979_ rbzero.wall_tracer.trackDistY\[-5\] vssd1 vssd1 vccd1 vccd1 _04989_
+ sky130_fd_sc_hd__nor2_1
XFILLER_141_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14034_ _06717_ _06718_ _06722_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__a21o_1
XFILLER_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18911_ rbzero.pov.spi_buffer\[5\] rbzero.pov.ready_buffer\[5\] _02608_ vssd1 vssd1
+ vccd1 vccd1 _02614_ sky130_fd_sc_hd__mux2_1
XFILLER_84_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11246_ _03941_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__clkbuf_4
XTAP_7051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19891_ _03111_ vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__clkinv_2
XTAP_7062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18842_ _02558_ _02559_ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__nor2_1
XTAP_7095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11177_ _03879_ _03894_ _03895_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__or3_4
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15985_ _08593_ _08597_ vssd1 vssd1 vccd1 vccd1 _08598_ sky130_fd_sc_hd__nand2_1
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18773_ _02492_ _02494_ _02166_ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__o21ai_1
XTAP_5660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17724_ _10030_ _10032_ _10031_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__o21ba_1
XTAP_5693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14936_ _07549_ vssd1 vssd1 vccd1 vccd1 _07550_ sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17655_ _10071_ _10079_ _01439_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__a21oi_1
X_14867_ _07478_ _07480_ _07349_ vssd1 vssd1 vccd1 vccd1 _07481_ sky130_fd_sc_hd__a21o_2
XFILLER_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16606_ _09063_ _09065_ vssd1 vssd1 vccd1 vccd1 _09215_ sky130_fd_sc_hd__and2_1
X_13818_ _06497_ _06506_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__nand2_1
X_17586_ _10118_ _10119_ _10121_ vssd1 vssd1 vccd1 vccd1 _10123_ sky130_fd_sc_hd__a21o_1
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14798_ rbzero.debug_overlay.playerX\[-5\] _07365_ rbzero.debug_overlay.playerX\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__o21ai_1
X_16537_ _09144_ _09145_ vssd1 vssd1 vccd1 vccd1 _09146_ sky130_fd_sc_hd__and2b_1
X_19325_ rbzero.pov.spi_counter\[6\] _02852_ _02854_ vssd1 vssd1 vccd1 vccd1 _00814_
+ sky130_fd_sc_hd__o21a_1
XFILLER_232_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13749_ _06435_ _06306_ _06437_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__o21ai_1
XFILLER_177_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16468_ _09075_ _09076_ _09034_ vssd1 vssd1 vccd1 vccd1 _09078_ sky130_fd_sc_hd__a21o_1
X_19256_ rbzero.spi_registers.got_new_leak _02742_ _02740_ _02811_ vssd1 vssd1 vccd1
+ vccd1 _00788_ sky130_fd_sc_hd__a31o_1
XFILLER_176_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18207_ _01923_ _01986_ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__xnor2_1
X_15419_ _08003_ _08031_ vssd1 vssd1 vccd1 vccd1 _08033_ sky130_fd_sc_hd__nor2_1
XFILLER_164_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19187_ _02771_ vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__clkbuf_1
X_16399_ _08994_ _09008_ vssd1 vssd1 vccd1 vccd1 _09009_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18138_ _01825_ _01917_ _01918_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__a21oi_1
XFILLER_145_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18069_ _01836_ _01749_ _01848_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__and3_1
XFILLER_208_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20100_ _03093_ _03135_ _03136_ _03137_ rbzero.texV\[-12\] vssd1 vssd1 vccd1 vccd1
+ _01306_ sky130_fd_sc_hd__a32o_1
XFILLER_99_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21080_ _00129_ _01096_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20031_ _03126_ vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__clkinv_2
XFILLER_8_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20933_ net69 _00949_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[70\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20864_ net79 _00880_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20795_ net84 _00811_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_224_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21347_ _00370_ _01363_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11100_ _03816_ _03817_ _03791_ _03819_ _00000_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__a41o_1
XFILLER_190_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12080_ net24 _04787_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__or2_1
XFILLER_172_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21278_ _00327_ _01294_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11031_ rbzero.map_rom.f4 _03733_ rbzero.map_rom.d6 rbzero.map_rom.f3 vssd1 vssd1
+ vccd1 vccd1 _03759_ sky130_fd_sc_hd__o2bb2a_1
X_20229_ rbzero.traced_texa\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _03245_
+ sky130_fd_sc_hd__or2_1
XFILLER_81_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15770_ _08357_ _08381_ vssd1 vssd1 vccd1 vccd1 _08384_ sky130_fd_sc_hd__and2_1
XFILLER_40_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12982_ _05471_ _05474_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__nand2_4
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14721_ _03800_ _07246_ _07335_ _07257_ vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__o211a_1
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11933_ net9 net10 vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__and2b_1
XFILLER_245_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _04939_ _09051_ _09610_ vssd1 vssd1 vccd1 vccd1 _09978_ sky130_fd_sc_hd__o21a_2
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ rbzero.wall_tracer.trackDistX\[7\] rbzero.wall_tracer.trackDistY\[7\] _05025_
+ vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__mux2_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11864_ rbzero.tex_b1\[5\] rbzero.tex_b1\[4\] _04544_ vssd1 vssd1 vccd1 vccd1 _04578_
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _06236_ _06246_ _06279_ _06280_ _06282_ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__a32o_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ _09901_ _09902_ _09908_ vssd1 vssd1 vccd1 vccd1 _09909_ sky130_fd_sc_hd__a21oi_1
XFILLER_220_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10815_ rbzero.tex_g0\[24\] rbzero.tex_g0\[23\] _03627_ vssd1 vssd1 vccd1 vccd1 _03632_
+ sky130_fd_sc_hd__mux2_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14583_ _03797_ _03778_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__and2_1
X_11795_ rbzero.tex_b0\[11\] _04142_ _04144_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__and3_1
XFILLER_60_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16322_ _08931_ _08932_ vssd1 vssd1 vccd1 vccd1 _08933_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19110_ rbzero.spi_registers.got_new_other _02721_ vssd1 vssd1 vccd1 vccd1 _02722_
+ sky130_fd_sc_hd__and2_1
XFILLER_213_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13534_ _05839_ _05878_ _06217_ vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__and3_1
XFILLER_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10746_ _03595_ vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19041_ rbzero.pov.spi_buffer\[67\] rbzero.pov.ready_buffer\[67\] _02673_ vssd1 vssd1
+ vccd1 vccd1 _02682_ sky130_fd_sc_hd__mux2_1
X_16253_ _08751_ _08753_ _08749_ vssd1 vssd1 vccd1 vccd1 _08864_ sky130_fd_sc_hd__a21bo_1
XFILLER_186_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13465_ _06152_ _06149_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__nor2_1
XFILLER_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10677_ _03559_ vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15204_ _07453_ rbzero.wall_tracer.stepDistY\[5\] vssd1 vssd1 vccd1 vccd1 _07818_
+ sky130_fd_sc_hd__nand2_1
XFILLER_127_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12416_ _05053_ _05056_ _05107_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__and3_1
XFILLER_51_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16184_ _08794_ _08795_ vssd1 vssd1 vccd1 vccd1 _08796_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13396_ _06083_ _06084_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15135_ _07442_ _07379_ _07399_ _07735_ vssd1 vssd1 vccd1 vccd1 _07749_ sky130_fd_sc_hd__or4_1
XFILLER_177_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12347_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__and2_1
XFILLER_86_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15066_ _07675_ vssd1 vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__clkbuf_4
XFILLER_142_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19943_ _03117_ vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__clkinv_2
X_12278_ _04965_ rbzero.wall_tracer.trackDistY\[-9\] _04966_ rbzero.wall_tracer.trackDistY\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__a22o_1
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14017_ _06696_ _06703_ _06705_ vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__a21oi_2
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11229_ _03868_ _03894_ _03897_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__or3_1
X_19874_ _03110_ vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__clkinv_2
XFILLER_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18825_ _02509_ rbzero.wall_tracer.rayAddendY\[8\] vssd1 vssd1 vccd1 vccd1 _02544_
+ sky130_fd_sc_hd__xor2_1
XTAP_6180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18756_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.debug_overlay.vplaneY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__and2_1
XTAP_5490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15968_ _08571_ _08572_ _08581_ vssd1 vssd1 vccd1 vccd1 _08582_ sky130_fd_sc_hd__o21ai_2
XFILLER_114_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17707_ _01488_ _01490_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__nand2_1
XFILLER_224_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14919_ rbzero.debug_overlay.playerY\[-3\] _07404_ vssd1 vssd1 vccd1 vccd1 _07533_
+ sky130_fd_sc_hd__nand2_1
X_15899_ _07442_ _07355_ _07552_ _07550_ vssd1 vssd1 vccd1 vccd1 _08513_ sky130_fd_sc_hd__or4_1
X_18687_ rbzero.wall_tracer.rayAddendY\[-2\] _00013_ _02412_ _02415_ vssd1 vssd1 vccd1
+ vccd1 _00615_ sky130_fd_sc_hd__o22a_1
XFILLER_188_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17638_ _09684_ _08723_ _10057_ _10059_ vssd1 vssd1 vccd1 vccd1 _10174_ sky130_fd_sc_hd__o31a_1
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17569_ _10103_ _10105_ vssd1 vssd1 vccd1 vccd1 _10106_ sky130_fd_sc_hd__xor2_1
XFILLER_210_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19308_ rbzero.pov.spi_counter\[2\] rbzero.pov.spi_counter\[1\] rbzero.pov.spi_counter\[0\]
+ _02842_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__and4bb_1
X_20580_ net88 _00596_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19239_ _02795_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__inv_2
XFILLER_108_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21201_ _00250_ _01217_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21132_ _00181_ _01148_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21063_ _00112_ _01079_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_232_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20014_ _03114_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__buf_4
XFILLER_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20916_ net69 _00932_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[53\] sky130_fd_sc_hd__dfxtp_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20847_ _00065_ _00863_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10600_ _03388_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__clkbuf_4
XFILLER_74_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11580_ _04108_ _04288_ _04297_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__and3_1
XFILLER_126_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20778_ net88 _00794_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout64 net72 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout75 net77 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout86 net89 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__buf_2
XFILLER_211_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout97 net98 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10531_ rbzero.tex_r0\[31\] rbzero.tex_r0\[30\] _03479_ vssd1 vssd1 vccd1 vccd1 _03483_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13250_ _05894_ _05897_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10462_ net48 rbzero.tex_r0\[63\] _03446_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__mux2_1
XFILLER_108_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12201_ net35 _04115_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__nand2_1
XFILLER_170_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13181_ _05775_ _05869_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__xor2_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10393_ _03408_ vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12132_ net30 _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__or2_1
XFILLER_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16940_ _09211_ _09212_ vssd1 vssd1 vccd1 vccd1 _09482_ sky130_fd_sc_hd__and2b_1
XFILLER_150_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12063_ _04768_ _04118_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__nor2_1
XFILLER_133_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11014_ rbzero.map_rom.f4 vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__inv_2
XFILLER_238_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16871_ _09404_ _09412_ vssd1 vssd1 vccd1 vccd1 _09413_ sky130_fd_sc_hd__xnor2_1
XFILLER_133_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18610_ _02346_ vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15822_ _08399_ _08405_ vssd1 vssd1 vccd1 vccd1 _08436_ sky130_fd_sc_hd__nand2_1
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19590_ rbzero.pov.ready_buffer\[63\] _07395_ _02962_ vssd1 vssd1 vccd1 vccd1 _02970_
+ sky130_fd_sc_hd__mux2_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15753_ _07880_ _07843_ _08366_ _08336_ vssd1 vssd1 vccd1 vccd1 _08367_ sky130_fd_sc_hd__o22a_1
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18541_ _02264_ _02269_ _02283_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__a21oi_1
XFILLER_246_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12965_ _05642_ _05653_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__nand2_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14704_ _07326_ vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11916_ _04625_ _04626_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__or2_1
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15684_ _07507_ _07879_ _07645_ _07718_ vssd1 vssd1 vccd1 vccd1 _08298_ sky130_fd_sc_hd__or4_1
X_18472_ _02203_ _02205_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__or2b_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _05487_ _05535_ _05578_ _05497_ _05584_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__a221o_1
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _07553_ _09055_ vssd1 vssd1 vccd1 vccd1 _09961_ sky130_fd_sc_hd__and2_1
X_14635_ rbzero.wall_tracer.trackDistX\[2\] rbzero.wall_tracer.trackDistY\[2\] _07258_
+ vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__mux2_1
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ rbzero.tex_b1\[27\] rbzero.tex_b1\[26\] _03934_ vssd1 vssd1 vccd1 vccd1 _04561_
+ sky130_fd_sc_hd__mux2_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14566_ rbzero.wall_tracer.stepDistY\[8\] _07234_ _04925_ vssd1 vssd1 vccd1 vccd1
+ _07235_ sky130_fd_sc_hd__mux2_1
X_17354_ _09889_ _09890_ _09891_ vssd1 vssd1 vccd1 vccd1 _09893_ sky130_fd_sc_hd__nand3_1
XFILLER_158_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11778_ rbzero.tex_b0\[21\] rbzero.tex_b0\[20\] _04001_ vssd1 vssd1 vccd1 vccd1 _04493_
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16305_ _07824_ _08793_ vssd1 vssd1 vccd1 vccd1 _08916_ sky130_fd_sc_hd__and2_1
XFILLER_207_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13517_ _06204_ _06205_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__and2_1
XFILLER_140_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17285_ _09791_ _09823_ vssd1 vssd1 vccd1 vccd1 _09824_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10729_ _03586_ vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__clkbuf_1
X_14497_ _07102_ _07179_ vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__nand2_2
XFILLER_144_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16236_ _08728_ _08743_ _08741_ vssd1 vssd1 vccd1 vccd1 _08847_ sky130_fd_sc_hd__a21o_1
XFILLER_174_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19024_ _02606_ vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__clkbuf_4
X_13448_ _05793_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__clkbuf_4
XFILLER_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16167_ _07814_ vssd1 vssd1 vccd1 vccd1 _08779_ sky130_fd_sc_hd__clkinv_2
XFILLER_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13379_ _06040_ _06054_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15118_ _07334_ _05078_ _07731_ _04932_ vssd1 vssd1 vccd1 vccd1 _07732_ sky130_fd_sc_hd__a211o_1
XFILLER_115_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16098_ _08459_ _08563_ _08697_ _08698_ _08709_ vssd1 vssd1 vccd1 vccd1 _08710_ sky130_fd_sc_hd__a41o_2
XFILLER_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15049_ _07661_ _07662_ vssd1 vssd1 vccd1 vccd1 _07663_ sky130_fd_sc_hd__nand2_4
XFILLER_142_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19926_ _03114_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__buf_4
XFILLER_69_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19857_ _03108_ vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__clkinv_2
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18808_ _02509_ rbzero.wall_tracer.rayAddendY\[7\] vssd1 vssd1 vccd1 vccd1 _02528_
+ sky130_fd_sc_hd__nand2_1
XFILLER_3_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19788_ _02753_ _02718_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__nor2_1
XFILLER_7_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18739_ _02462_ _02460_ _02461_ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__and3_1
XFILLER_92_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20701_ net87 _00717_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20632_ net55 _00648_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20563_ net136 _00579_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20494_ net111 _00510_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21115_ _00164_ _01131_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_6938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21046_ _00095_ _01062_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12750_ _05417_ _05438_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__nor2_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _04007_ _04412_ _04416_ _03956_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__a211o_1
XFILLER_42_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12681_ _03790_ _05242_ _05244_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__a21o_2
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _05517_ _07107_ _07108_ vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__and3_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11632_ rbzero.tex_g0\[59\] _04142_ _04144_ _03929_ vssd1 vssd1 vccd1 vccd1 _04349_
+ sky130_fd_sc_hd__a31o_1
XFILLER_168_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14351_ _05431_ _07020_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__nand2_1
XFILLER_50_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11563_ rbzero.debug_overlay.playerY\[-4\] _04242_ _04238_ rbzero.debug_overlay.playerY\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__a22o_1
XFILLER_11_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13302_ _05884_ _05990_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__and2_1
X_17070_ _04939_ _09051_ _09610_ vssd1 vssd1 vccd1 vccd1 _09611_ sky130_fd_sc_hd__o21ai_4
XFILLER_196_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10514_ rbzero.tex_r0\[39\] rbzero.tex_r0\[38\] _03468_ vssd1 vssd1 vccd1 vccd1 _03474_
+ sky130_fd_sc_hd__mux2_1
X_14282_ _06631_ _06689_ vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__or2b_1
XFILLER_183_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11494_ _04199_ _04210_ _04211_ _04196_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__or4b_1
X_16021_ _04929_ _08633_ vssd1 vssd1 vccd1 vccd1 _08634_ sky130_fd_sc_hd__nand2_4
XFILLER_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13233_ _05909_ _05921_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10445_ rbzero.tex_r1\[5\] rbzero.tex_r1\[6\] _03433_ vssd1 vssd1 vccd1 vccd1 _03436_
+ sky130_fd_sc_hd__mux2_1
XFILLER_237_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13164_ _05739_ _05852_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10376_ _03399_ vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__clkbuf_1
X_12115_ _04820_ o_rgb[14] _04821_ net31 vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__o211a_1
XFILLER_237_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17972_ _01733_ _01753_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__xnor2_1
X_13095_ _05781_ _05783_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__xor2_1
XFILLER_215_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19711_ _02708_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__buf_4
X_16923_ _09464_ vssd1 vssd1 vccd1 vccd1 _09465_ sky130_fd_sc_hd__clkbuf_2
XFILLER_133_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12046_ net4 net3 vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__and2b_1
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19642_ _03009_ _03008_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__nand2_1
XFILLER_238_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16854_ _09394_ _09395_ vssd1 vssd1 vccd1 vccd1 _09396_ sky130_fd_sc_hd__xor2_1
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15805_ _07517_ _08394_ _07842_ _08395_ vssd1 vssd1 vccd1 vccd1 _08419_ sky130_fd_sc_hd__or4b_1
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19573_ rbzero.debug_overlay.playerX\[-9\] vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__inv_2
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13997_ _06632_ _06685_ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__or2_1
X_16785_ rbzero.wall_tracer.trackDistX\[-5\] rbzero.wall_tracer.stepDistX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _09332_ sky130_fd_sc_hd__or2_1
XFILLER_4_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18524_ _02260_ _02267_ _02265_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__a21o_1
XFILLER_98_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15736_ _08330_ _08348_ _08349_ vssd1 vssd1 vccd1 vccd1 _08350_ sky130_fd_sc_hd__a21oi_1
X_12948_ _05634_ _05636_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__and2_1
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18455_ rbzero.debug_overlay.vplaneX\[0\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__or2_1
XFILLER_221_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15667_ _08278_ _08279_ vssd1 vssd1 vccd1 vccd1 _08281_ sky130_fd_sc_hd__or2_1
X_12879_ _05440_ _05405_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__nor2_2
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17406_ _09932_ _09943_ vssd1 vssd1 vccd1 vccd1 _09944_ sky130_fd_sc_hd__nand2_1
XFILLER_222_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14618_ _07245_ _07273_ _07274_ _07251_ vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__o211a_1
XFILLER_61_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15598_ _08192_ _08211_ vssd1 vssd1 vccd1 vccd1 _08212_ sky130_fd_sc_hd__xnor2_1
X_18386_ rbzero.spi_registers.spi_done _03292_ _02140_ vssd1 vssd1 vccd1 vccd1 _02141_
+ sky130_fd_sc_hd__and3_1
XFILLER_226_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17337_ _09697_ _09747_ _09875_ vssd1 vssd1 vccd1 vccd1 _09876_ sky130_fd_sc_hd__a21oi_1
X_14549_ _07101_ _07220_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__nand2_1
XFILLER_193_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17268_ _09796_ _09806_ vssd1 vssd1 vccd1 vccd1 _09807_ sky130_fd_sc_hd__xor2_1
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19007_ _02664_ vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16219_ _08828_ _08830_ vssd1 vssd1 vccd1 vccd1 _08831_ sky130_fd_sc_hd__nor2_1
X_17199_ _09737_ _09738_ vssd1 vssd1 vccd1 vccd1 _09739_ sky130_fd_sc_hd__xor2_1
XFILLER_220_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19909_ _03113_ vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__clkinv_2
XFILLER_229_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20615_ net84 _00631_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20546_ net125 _00562_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20477_ net96 _00493_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10230_ rbzero.tex_b1\[43\] rbzero.tex_b1\[44\] _03322_ vssd1 vssd1 vccd1 vccd1 _03323_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13920_ _06608_ _06588_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21029_ net109 _01045_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_134_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13851_ _06168_ _06172_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__or2_1
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12802_ _05422_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__clkinv_2
XFILLER_74_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16570_ _09161_ _09178_ vssd1 vssd1 vccd1 vccd1 _09179_ sky130_fd_sc_hd__and2_1
X_13782_ _06260_ _06289_ _06303_ _06101_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__a211o_1
XFILLER_222_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10994_ _03725_ vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15521_ _07350_ _07353_ vssd1 vssd1 vccd1 vccd1 _08135_ sky130_fd_sc_hd__nand2_4
X_12733_ _05331_ _05332_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__or2_2
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15452_ _08058_ _08065_ vssd1 vssd1 vccd1 vccd1 _08066_ sky130_fd_sc_hd__xnor2_1
X_18240_ rbzero.wall_tracer.trackDistY\[-9\] rbzero.wall_tracer.stepDistY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__nand2_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12664_ _05339_ _05352_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__xnor2_4
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14403_ _06990_ _07053_ _07054_ _07091_ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__a31o_1
XFILLER_141_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11615_ rbzero.tex_g0\[11\] _04142_ _04144_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__and3_1
X_18171_ _07818_ _07823_ _08718_ vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__a21o_1
X_15383_ _07994_ _07996_ vssd1 vssd1 vccd1 vccd1 _07997_ sky130_fd_sc_hd__nand2_1
XFILLER_169_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12595_ _05220_ _05283_ _05280_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__a21o_1
XFILLER_15_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17122_ _09568_ _09587_ _09586_ vssd1 vssd1 vccd1 vccd1 _09662_ sky130_fd_sc_hd__a21o_1
XFILLER_204_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14334_ _07016_ _07022_ _06985_ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__mux2_1
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11546_ rbzero.debug_overlay.vplaneY\[-5\] _04214_ _04237_ rbzero.debug_overlay.vplaneY\[-6\]
+ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__a22o_1
XFILLER_102_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17053_ _09449_ _09451_ _09593_ vssd1 vssd1 vccd1 vccd1 _09594_ sky130_fd_sc_hd__o21ai_1
X_14265_ _06931_ _06943_ _06952_ _06953_ vssd1 vssd1 vccd1 vccd1 _06954_ sky130_fd_sc_hd__a211o_1
XFILLER_143_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11477_ gpout0.hpos\[3\] _03804_ gpout0.hpos\[4\] vssd1 vssd1 vccd1 vccd1 _04195_
+ sky130_fd_sc_hd__a21oi_1
X_16004_ _07472_ _07641_ _07400_ vssd1 vssd1 vccd1 vccd1 _08617_ sky130_fd_sc_hd__a21oi_2
X_13216_ _05817_ _05830_ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10428_ rbzero.tex_r1\[13\] rbzero.tex_r1\[14\] _03422_ vssd1 vssd1 vccd1 vccd1 _03427_
+ sky130_fd_sc_hd__mux2_1
X_14196_ _06310_ _06634_ _06884_ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__or3_1
XFILLER_171_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13147_ _05825_ _05829_ _05835_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__o21a_1
XFILLER_124_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ rbzero.tex_r1\[46\] rbzero.tex_r1\[47\] _03389_ vssd1 vssd1 vccd1 vccd1 _03391_
+ sky130_fd_sc_hd__mux2_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ _08594_ _09603_ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__nor2_1
X_13078_ _05726_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__buf_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16906_ _08771_ _08788_ _09191_ _09447_ vssd1 vssd1 vccd1 vccd1 _09448_ sky130_fd_sc_hd__a31o_1
X_12029_ _04718_ net6 _04732_ _04734_ _04737_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__a32o_1
XFILLER_113_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17886_ _01551_ _01553_ _01550_ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__a21bo_1
XFILLER_152_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19625_ rbzero.pov.ready_buffer\[71\] _02963_ _02981_ _02996_ vssd1 vssd1 vccd1 vccd1
+ _02997_ sky130_fd_sc_hd__o211a_1
XFILLER_54_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16837_ _09156_ _09372_ _09378_ vssd1 vssd1 vccd1 vccd1 _09379_ sky130_fd_sc_hd__a21oi_1
XFILLER_113_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19556_ net52 rbzero.pov.mosi_buffer\[0\] _02708_ vssd1 vssd1 vccd1 vccd1 _02947_
+ sky130_fd_sc_hd__mux2_1
X_16768_ _07332_ _08571_ vssd1 vssd1 vccd1 vccd1 _09317_ sky130_fd_sc_hd__and2_1
XFILLER_206_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18507_ _02223_ _02239_ _02241_ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a21oi_1
XFILLER_202_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15719_ _08298_ _08294_ _08297_ vssd1 vssd1 vccd1 vccd1 _08333_ sky130_fd_sc_hd__nand3_1
XFILLER_179_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19487_ _02911_ vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__clkbuf_1
X_16699_ rbzero.traced_texa\[1\] _09264_ _09265_ rbzero.wall_tracer.visualWallDist\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__a22o_1
XFILLER_224_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18438_ _02166_ _02187_ _02188_ _09254_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a31o_1
XFILLER_167_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18369_ _02119_ _02122_ _02120_ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__o21ai_1
XFILLER_33_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20400_ net123 _00431_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21380_ net127 _01396_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20331_ _02727_ _03264_ _03265_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__and3_1
XFILLER_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20262_ _03255_ vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__clkinv_2
XFILLER_66_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20193_ _09245_ _03214_ _03215_ _03064_ rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1
+ _01321_ sky130_fd_sc_hd__a32o_1
XFILLER_130_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11400_ _04118_ vssd1 vssd1 vccd1 vccd1 o_rgb[6] sky130_fd_sc_hd__inv_2
X_12380_ _05071_ _05072_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__and2b_1
XFILLER_138_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11331_ _04048_ _04049_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__and2_1
X_20529_ net120 _00545_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14050_ _06699_ _06701_ vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__xor2_1
XFILLER_153_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11262_ rbzero.tex_r0\[34\] _03980_ _03942_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__a21o_1
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13001_ _05620_ _05689_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__and2_1
XFILLER_49_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10213_ rbzero.tex_b1\[51\] rbzero.tex_b1\[52\] _03311_ vssd1 vssd1 vccd1 vccd1 _03314_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11193_ rbzero.tex_r0\[55\] rbzero.tex_r0\[54\] _03904_ vssd1 vssd1 vccd1 vccd1 _03912_
+ sky130_fd_sc_hd__mux2_1
XTAP_6521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17740_ _10155_ _01523_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__xnor2_1
XFILLER_216_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14952_ _07560_ _07561_ _07565_ _04937_ vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__a22o_1
XFILLER_248_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13903_ _06530_ _06591_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__and2_1
X_17671_ _07886_ _10095_ _01454_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14883_ rbzero.debug_overlay.playerY\[-3\] _07404_ vssd1 vssd1 vccd1 vccd1 _07497_
+ sky130_fd_sc_hd__or2_1
XFILLER_235_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19410_ rbzero.pov.spi_buffer\[3\] rbzero.pov.spi_buffer\[4\] _02866_ vssd1 vssd1
+ vccd1 vccd1 _02871_ sky130_fd_sc_hd__mux2_1
XFILLER_235_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16622_ _08844_ _09094_ _09230_ vssd1 vssd1 vccd1 vccd1 _09231_ sky130_fd_sc_hd__a21o_1
X_13834_ _06462_ _06464_ _06463_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__a21o_1
XFILLER_169_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19341_ _02857_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__clkinv_2
X_16553_ _09035_ _09044_ _09043_ vssd1 vssd1 vccd1 vccd1 _09162_ sky130_fd_sc_hd__a21bo_1
X_13765_ _06450_ _06452_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__or2_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10977_ rbzero.tex_b0\[11\] rbzero.tex_b0\[10\] _03715_ vssd1 vssd1 vccd1 vccd1 _03717_
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15504_ _07378_ _07399_ _07508_ _07575_ vssd1 vssd1 vccd1 vccd1 _08118_ sky130_fd_sc_hd__nor4_1
XFILLER_71_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12716_ _05399_ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__nor2_2
X_19272_ _02820_ vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__clkbuf_1
XFILLER_245_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16484_ _09091_ _09093_ vssd1 vssd1 vccd1 vccd1 _09094_ sky130_fd_sc_hd__xnor2_1
X_13696_ _06344_ _06346_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__xnor2_2
XFILLER_188_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18223_ _01997_ _01998_ _01999_ _02001_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__a31o_1
XFILLER_176_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15435_ _07377_ _07485_ _07574_ _07398_ vssd1 vssd1 vccd1 vccd1 _08049_ sky130_fd_sc_hd__o22a_1
X_12647_ _05233_ _05263_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__or2_2
XFILLER_203_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18154_ _01736_ _01847_ _01849_ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__a21oi_1
XFILLER_175_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15366_ _07968_ _07978_ _07979_ vssd1 vssd1 vccd1 vccd1 _07980_ sky130_fd_sc_hd__a21bo_1
XFILLER_89_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12578_ _05266_ _05172_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__xnor2_2
XFILLER_106_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17105_ _09642_ _09643_ _09644_ vssd1 vssd1 vccd1 vccd1 _09646_ sky130_fd_sc_hd__and3_1
XFILLER_157_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14317_ _06990_ _07005_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__nand2_1
XFILLER_157_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11529_ rbzero.debug_overlay.facingX\[-2\] _04245_ _04103_ _04246_ vssd1 vssd1 vccd1
+ vccd1 _04247_ sky130_fd_sc_hd__a211o_1
X_15297_ _07910_ vssd1 vssd1 vccd1 vccd1 _07911_ sky130_fd_sc_hd__inv_2
X_18085_ _01767_ _01768_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__nand2_1
XFILLER_176_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17036_ _07696_ _08640_ _07890_ vssd1 vssd1 vccd1 vccd1 _09577_ sky130_fd_sc_hd__a21oi_2
X_14248_ _06935_ _06936_ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__xor2_1
XFILLER_217_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14179_ _06857_ _06863_ _06867_ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__o21a_1
XFILLER_113_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ rbzero.pov.spi_buffer\[41\] rbzero.pov.ready_buffer\[41\] _02651_ vssd1 vssd1
+ vccd1 vccd1 _02654_ sky130_fd_sc_hd__mux2_1
XFILLER_140_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17938_ _03797_ _01719_ _01720_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__or3b_2
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17869_ _09429_ _08852_ _01529_ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__o21ba_1
XFILLER_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19608_ rbzero.debug_overlay.playerX\[0\] _07562_ vssd1 vssd1 vccd1 vccd1 _02983_
+ sky130_fd_sc_hd__nand2_1
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20880_ net58 _00896_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19539_ _02938_ vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__clkbuf_1
XFILLER_241_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21363_ _00386_ _01379_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20314_ rbzero.traced_texVinit\[4\] _09266_ _03259_ _09261_ vssd1 vssd1 vccd1 vccd1
+ _01398_ sky130_fd_sc_hd__a22o_1
XFILLER_135_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21294_ net134 _01310_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20245_ _03253_ vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__clkinv_2
XFILLER_104_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20176_ _03194_ _03198_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__nand2_1
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10900_ _03676_ vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__clkbuf_1
XFILLER_217_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11880_ _04592_ _03289_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__nand2_1
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10831_ _03640_ vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13550_ _05433_ _05608_ _05611_ _05583_ vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__or4_1
XFILLER_242_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10762_ _03603_ vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12501_ _05189_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__buf_2
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13481_ _06150_ _06153_ _06148_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10693_ rbzero.tex_g1\[17\] rbzero.tex_g1\[18\] _03563_ vssd1 vssd1 vccd1 vccd1 _03568_
+ sky130_fd_sc_hd__mux2_1
XFILLER_197_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15220_ _04928_ _07832_ _07651_ _07833_ vssd1 vssd1 vccd1 vccd1 _07834_ sky130_fd_sc_hd__a31oi_4
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12432_ _05122_ _05123_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__and2_1
XFILLER_205_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15151_ _07470_ _07735_ vssd1 vssd1 vccd1 vccd1 _07765_ sky130_fd_sc_hd__nor2_1
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12363_ _05048_ _05052_ _05055_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__o21ai_2
XFILLER_103_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14102_ _06786_ _06790_ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__and2_1
XFILLER_165_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11314_ rbzero.floor_leak\[1\] _03914_ _04032_ rbzero.floor_leak\[0\] vssd1 vssd1
+ vccd1 vccd1 _04033_ sky130_fd_sc_hd__o211a_1
X_15082_ _07686_ _07695_ _04928_ vssd1 vssd1 vccd1 vccd1 _07696_ sky130_fd_sc_hd__o21ai_4
XFILLER_114_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12294_ _04984_ _04987_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__or2_1
XFILLER_154_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14033_ _05668_ _06321_ _06720_ _06721_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__a31o_1
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18910_ _02613_ vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__clkbuf_1
XTAP_7030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11245_ _03939_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__buf_2
XTAP_7041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19890_ _03111_ vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__clkinv_2
XFILLER_107_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18841_ _02557_ _02555_ _02556_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__nor3_1
XTAP_7085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ _03834_ _03872_ _03878_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__nor3b_2
XTAP_6351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18772_ _02492_ _02494_ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__and2_1
XTAP_6395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15984_ _07388_ _08594_ _08595_ _08596_ vssd1 vssd1 vccd1 vccd1 _08597_ sky130_fd_sc_hd__o22ai_1
XTAP_5650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17723_ rbzero.wall_tracer.trackDistX\[6\] rbzero.wall_tracer.stepDistX\[6\] vssd1
+ vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__and2_1
XFILLER_208_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14935_ _04936_ _07545_ _07548_ vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__o21ai_2
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17654_ _10078_ _10072_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__and2b_1
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14866_ _07346_ _07479_ vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__nand2_1
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16605_ _09206_ _09213_ vssd1 vssd1 vccd1 vccd1 _09214_ sky130_fd_sc_hd__xnor2_1
XFILLER_224_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13817_ _06495_ _06496_ vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__or2_1
X_17585_ _10118_ _10119_ _10121_ vssd1 vssd1 vccd1 vccd1 _10122_ sky130_fd_sc_hd__nand3_1
X_14797_ rbzero.debug_overlay.playerX\[-4\] rbzero.debug_overlay.playerX\[-5\] _07365_
+ vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__or3_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19324_ rbzero.pov.spi_counter\[6\] _02852_ _02844_ vssd1 vssd1 vccd1 vccd1 _02854_
+ sky130_fd_sc_hd__a21boi_1
X_16536_ _08086_ _08223_ _07597_ _07620_ vssd1 vssd1 vccd1 vccd1 _09145_ sky130_fd_sc_hd__or4_1
X_13748_ _06380_ _06436_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__or2_1
XFILLER_56_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19255_ _02804_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__inv_2
X_16467_ _09034_ _09075_ _09076_ vssd1 vssd1 vccd1 vccd1 _09077_ sky130_fd_sc_hd__nand3_1
X_13679_ _05434_ _06307_ _06308_ _06367_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__nor4_4
XFILLER_32_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18206_ _01924_ _01985_ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15418_ _08003_ _08031_ vssd1 vssd1 vccd1 vccd1 _08032_ sky130_fd_sc_hd__xor2_1
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19186_ _09247_ _02770_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__and2_1
X_16398_ _09006_ _09007_ vssd1 vssd1 vccd1 vccd1 _09008_ sky130_fd_sc_hd__nor2_1
XFILLER_191_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18137_ rbzero.wall_tracer.trackDistX\[10\] rbzero.wall_tracer.stepDistX\[10\] vssd1
+ vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15349_ _07604_ _07962_ vssd1 vssd1 vccd1 vccd1 _07963_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18068_ _01836_ _01749_ _01848_ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a21oi_1
XFILLER_172_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17019_ _09556_ _09558_ vssd1 vssd1 vccd1 vccd1 _09560_ sky130_fd_sc_hd__and2_1
XFILLER_176_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20030_ _03126_ vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__clkinv_2
XFILLER_217_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20932_ net67 _00948_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[69\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20863_ net79 _00879_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20794_ net84 _00810_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21346_ _00369_ _01362_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21277_ _00326_ _01293_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11030_ rbzero.map_rom.f1 rbzero.map_rom.c6 vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__nand2_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20228_ _09245_ _03243_ _03244_ _03064_ rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1
+ _01327_ sky130_fd_sc_hd__a32o_1
XFILLER_231_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20159_ rbzero.texV\[-2\] _02989_ _03142_ _03186_ vssd1 vssd1 vccd1 vccd1 _01316_
+ sky130_fd_sc_hd__a22o_1
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _05668_ _05669_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__xnor2_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14720_ _07334_ _03799_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__nand2_1
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11932_ net10 net9 vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__and2b_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14651_ _03800_ _07296_ _07297_ _07257_ vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__o211a_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ _03920_ _04572_ _04576_ _03949_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__a211o_1
XFILLER_79_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13602_ _06283_ _06265_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__and2b_1
X_10814_ _03631_ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__clkbuf_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _09906_ _09907_ vssd1 vssd1 vccd1 vccd1 _09908_ sky130_fd_sc_hd__nand2_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14582_ rbzero.wall_tracer.trackDistX\[-12\] rbzero.wall_tracer.trackDistY\[-12\]
+ _07246_ vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__mux2_1
X_11794_ rbzero.tex_b0\[9\] rbzero.tex_b0\[8\] _03925_ vssd1 vssd1 vccd1 vccd1 _04509_
+ sky130_fd_sc_hd__mux2_1
XFILLER_232_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16321_ _07847_ _08787_ vssd1 vssd1 vccd1 vccd1 _08932_ sky130_fd_sc_hd__nor2_1
XFILLER_242_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13533_ _06176_ _06221_ vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__or2_2
X_10745_ rbzero.tex_g0\[57\] rbzero.tex_g0\[56\] _03593_ vssd1 vssd1 vccd1 vccd1 _03595_
+ sky130_fd_sc_hd__mux2_1
XFILLER_199_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19040_ _02681_ vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16252_ _08733_ _08736_ _08731_ vssd1 vssd1 vccd1 vccd1 _08863_ sky130_fd_sc_hd__a21bo_1
X_13464_ _06151_ _06149_ _06152_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__a21o_1
X_10676_ rbzero.tex_g1\[25\] rbzero.tex_g1\[26\] _03552_ vssd1 vssd1 vccd1 vccd1 _03559_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15203_ _07816_ vssd1 vssd1 vccd1 vccd1 _07817_ sky130_fd_sc_hd__clkbuf_4
X_12415_ _05053_ _05056_ _05107_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16183_ _08335_ _08645_ vssd1 vssd1 vccd1 vccd1 _08795_ sky130_fd_sc_hd__nor2_1
X_13395_ _06032_ _06034_ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15134_ _07379_ _07736_ vssd1 vssd1 vccd1 vccd1 _07748_ sky130_fd_sc_hd__nor2_1
X_12346_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__xor2_2
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15065_ _07678_ _07664_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__nor2_1
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19942_ _03117_ vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__clkinv_2
X_12277_ _04968_ rbzero.wall_tracer.trackDistY\[-11\] _04970_ vssd1 vssd1 vccd1 vccd1
+ _04971_ sky130_fd_sc_hd__a21o_1
XFILLER_218_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14016_ _06639_ _06704_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__nand2_1
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11228_ _03932_ _03933_ _03937_ _03943_ _03946_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__o221a_1
XFILLER_214_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19873_ _03110_ vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__clkinv_2
XFILLER_218_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18824_ rbzero.wall_tracer.rayAddendY\[7\] _00013_ _02543_ vssd1 vssd1 vccd1 vccd1
+ _00624_ sky130_fd_sc_hd__o21a_1
XFILLER_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11159_ _03876_ _03877_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18755_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.debug_overlay.vplaneY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__nor2_1
XTAP_5480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15967_ _08571_ _08572_ _08579_ _08580_ vssd1 vssd1 vccd1 vccd1 _08581_ sky130_fd_sc_hd__a211o_1
XFILLER_49_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17706_ _01488_ _01490_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__nor2_1
XFILLER_208_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14918_ _07530_ _07531_ vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__and2_1
XFILLER_209_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18686_ _02166_ _02413_ _02414_ _09254_ vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__a31o_1
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15898_ _08509_ _08511_ vssd1 vssd1 vccd1 vccd1 _08512_ sky130_fd_sc_hd__xnor2_2
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17637_ _10171_ _10172_ vssd1 vssd1 vccd1 vccd1 _10173_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14849_ rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\] rbzero.debug_overlay.playerX\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__o21ai_1
XFILLER_149_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17568_ _09968_ _08917_ _09965_ _10104_ vssd1 vssd1 vccd1 vccd1 _10105_ sky130_fd_sc_hd__o31a_1
XFILLER_205_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19307_ rbzero.pov.spi_counter\[5\] rbzero.pov.spi_counter\[4\] rbzero.pov.spi_counter\[3\]
+ rbzero.pov.spi_counter\[6\] vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__and4bb_1
X_16519_ _09126_ _09127_ vssd1 vssd1 vccd1 vccd1 _09128_ sky130_fd_sc_hd__xnor2_1
XFILLER_210_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17499_ _10011_ _10013_ vssd1 vssd1 vccd1 vccd1 _10036_ sky130_fd_sc_hd__or2_1
XFILLER_149_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19238_ _02801_ vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__clkbuf_1
XFILLER_149_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19169_ rbzero.spi_registers.new_sky\[4\] rbzero.spi_registers.got_new_sky _02724_
+ _02753_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__a31o_1
XFILLER_129_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21200_ _00249_ _01216_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21131_ _00180_ _01147_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21062_ _00111_ _01078_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20013_ _03123_ vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__clkinv_2
XFILLER_87_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20915_ net68 _00931_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[52\] sky130_fd_sc_hd__dfxtp_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20846_ _00064_ _00862_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout54 net59 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_2
X_20777_ net102 _00793_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout65 net72 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout76 net77 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10530_ _03482_ vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout87 net88 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_2
XFILLER_122_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout98 net141 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_4
XFILLER_202_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10461_ _03445_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__clkbuf_4
XFILLER_136_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12200_ _04872_ _04903_ _04905_ _04885_ _04895_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__a221o_1
XFILLER_108_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13180_ _05858_ _05868_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10392_ rbzero.tex_r1\[30\] rbzero.tex_r1\[31\] _03400_ vssd1 vssd1 vccd1 vccd1 _03408_
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12131_ _03294_ _03295_ gpout0.vpos\[8\] _04110_ net27 _04832_ vssd1 vssd1 vccd1
+ vccd1 _04838_ sky130_fd_sc_hd__mux4_1
X_21329_ _00352_ _01345_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12062_ _04768_ o_rgb[14] _04769_ net25 vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__o211a_1
XFILLER_78_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11013_ rbzero.map_rom.f3 rbzero.map_rom.c6 vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__nand2_1
XFILLER_46_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16870_ _09406_ _09411_ vssd1 vssd1 vccd1 vccd1 _09412_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15821_ _08418_ _08424_ _08427_ _08434_ _08406_ vssd1 vssd1 vccd1 vccd1 _08435_ sky130_fd_sc_hd__a221o_1
XFILLER_133_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18540_ _02264_ _02269_ _02283_ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__and3_1
X_15752_ _07789_ _07593_ _07838_ _08293_ vssd1 vssd1 vccd1 vccd1 _08366_ sky130_fd_sc_hd__and4bb_1
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _05651_ _05652_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__or2_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14703_ rbzero.wall_tracer.stepDistX\[6\] _07225_ _07316_ vssd1 vssd1 vccd1 vccd1
+ _07326_ sky130_fd_sc_hd__mux2_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ _04078_ _03781_ _03784_ _03291_ net9 _04618_ vssd1 vssd1 vccd1 vccd1 _04626_
+ sky130_fd_sc_hd__mux4_1
X_18471_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__or2_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15683_ _08296_ _07842_ vssd1 vssd1 vccd1 vccd1 _08297_ sky130_fd_sc_hd__nor2_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _05497_ _05496_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__nor2_1
XFILLER_2_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17422_ _09958_ _09959_ vssd1 vssd1 vccd1 vccd1 _09960_ sky130_fd_sc_hd__xnor2_1
XFILLER_205_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14634_ _07245_ _07284_ _07285_ _07251_ vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__o211a_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _04556_ _04559_ _03920_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__mux2_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17353_ _09889_ _09890_ _09891_ vssd1 vssd1 vccd1 vccd1 _09892_ sky130_fd_sc_hd__a21o_1
XFILLER_183_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ _07098_ _07233_ _07133_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__a21oi_4
X_11777_ _04490_ _04491_ _03968_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__mux2_1
XFILLER_198_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16304_ _08779_ _08788_ vssd1 vssd1 vccd1 vccd1 _08915_ sky130_fd_sc_hd__nand2_1
XFILLER_202_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13516_ _06196_ _06197_ _06203_ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__or3_1
XFILLER_119_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10728_ rbzero.tex_g1\[0\] rbzero.tex_g1\[1\] _03299_ vssd1 vssd1 vccd1 vccd1 _03586_
+ sky130_fd_sc_hd__mux2_1
X_17284_ _09807_ _09822_ vssd1 vssd1 vccd1 vccd1 _09823_ sky130_fd_sc_hd__xor2_1
X_14496_ _07174_ _07026_ _07175_ _07178_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_140_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19023_ _02672_ vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__clkbuf_1
X_16235_ _08844_ _08845_ vssd1 vssd1 vccd1 vccd1 _08846_ sky130_fd_sc_hd__nor2_1
XFILLER_220_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13447_ _06126_ _06134_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__nor2_1
X_10659_ rbzero.tex_g1\[33\] rbzero.tex_g1\[34\] _03541_ vssd1 vssd1 vccd1 vccd1 _03550_
+ sky130_fd_sc_hd__mux2_1
X_16166_ _08769_ _08777_ vssd1 vssd1 vccd1 vccd1 _08778_ sky130_fd_sc_hd__xor2_1
XFILLER_220_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13378_ _06064_ _06060_ _06063_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__and3_1
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15117_ _07334_ _05210_ vssd1 vssd1 vccd1 vccd1 _07731_ sky130_fd_sc_hd__nor2_1
XFILLER_177_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12329_ _04980_ _04964_ _04972_ _05022_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__or4_1
XFILLER_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16097_ _08589_ _08561_ _08696_ vssd1 vssd1 vccd1 vccd1 _08709_ sky130_fd_sc_hd__a21oi_1
XFILLER_173_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15048_ _03795_ rbzero.wall_tracer.stepDistY\[3\] _04928_ vssd1 vssd1 vccd1 vccd1
+ _07662_ sky130_fd_sc_hd__o21a_1
XFILLER_69_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19925_ _03115_ vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__clkinv_2
XFILLER_190_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19856_ _03108_ vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__clkinv_2
XFILLER_190_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18807_ _02287_ _02518_ _02519_ _02527_ vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__a31o_1
X_19787_ _04101_ _02716_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__or2_1
X_16999_ _09538_ _09539_ vssd1 vssd1 vccd1 vccd1 _09540_ sky130_fd_sc_hd__xor2_1
XFILLER_62_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18738_ _02460_ _02461_ _02462_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__a21oi_1
XFILLER_225_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18669_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.wall_tracer.rayAddendY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__nand2_1
XFILLER_93_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20700_ net87 _00716_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20631_ net55 _00647_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20562_ net136 _00578_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20493_ net111 _00509_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21114_ _00163_ _01130_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_6917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21045_ _00094_ _01061_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _03958_ _04413_ _04414_ _04415_ _03994_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__o221a_1
XFILLER_243_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12680_ _05365_ _05366_ _05367_ _05368_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__o22ai_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11631_ rbzero.tex_g0\[58\] _03974_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__and2_1
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20829_ _00047_ _00845_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14350_ _05593_ _07014_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__and2_1
XFILLER_168_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11562_ rbzero.debug_overlay.playerY\[-8\] _04218_ _04278_ rbzero.debug_overlay.playerY\[4\]
+ _04279_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__a221o_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13301_ _05793_ _05728_ _05819_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__o21ai_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10513_ _03473_ vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__clkbuf_1
X_14281_ _06794_ _06966_ _06969_ _06968_ vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__a31o_1
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11493_ _03290_ _03823_ _04204_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__a21boi_1
X_16020_ _08629_ rbzero.wall_tracer.stepDistY\[7\] _07694_ _08632_ vssd1 vssd1 vccd1
+ vccd1 _08633_ sky130_fd_sc_hd__a22o_4
XFILLER_183_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13232_ _05917_ _05920_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__nor2_1
XFILLER_104_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10444_ _03435_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13163_ _05847_ _05851_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10375_ rbzero.tex_r1\[38\] rbzero.tex_r1\[39\] _03389_ vssd1 vssd1 vccd1 vccd1 _03399_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12114_ _04820_ _04447_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__nand2_1
XFILLER_87_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17971_ _01735_ _01752_ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__xnor2_1
X_13094_ _05719_ _05734_ _05782_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__o21a_1
XFILLER_124_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19710_ _03062_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__buf_2
X_16922_ _07470_ _07971_ _09200_ vssd1 vssd1 vccd1 vccd1 _09464_ sky130_fd_sc_hd__or3_1
X_12045_ _04115_ _04753_ _04720_ gpout0.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _04754_
+ sky130_fd_sc_hd__a22o_1
XFILLER_238_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19641_ _03009_ rbzero.pov.ready_buffer\[44\] _02835_ vssd1 vssd1 vccd1 vccd1 _03010_
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16853_ _08510_ _08722_ vssd1 vssd1 vccd1 vccd1 _09395_ sky130_fd_sc_hd__nor2_1
XFILLER_78_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15804_ _08397_ _08401_ vssd1 vssd1 vccd1 vccd1 _08418_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19572_ _02955_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__clkbuf_4
X_16784_ _09279_ _08700_ vssd1 vssd1 vccd1 vccd1 _09331_ sky130_fd_sc_hd__nor2_1
XFILLER_207_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13996_ _06633_ _06680_ _06684_ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__o21a_1
XFILLER_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18523_ _02260_ _02265_ _02267_ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__and3_1
X_15735_ _08331_ _08347_ vssd1 vssd1 vccd1 vccd1 _08349_ sky130_fd_sc_hd__and2b_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ _05613_ _05635_ _05537_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__o21ai_4
XFILLER_65_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18454_ _02192_ _02195_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__nand2_1
X_15666_ _08278_ _08279_ vssd1 vssd1 vccd1 vccd1 _08280_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__buf_2
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17405_ _09941_ _09942_ vssd1 vssd1 vccd1 vccd1 _09943_ sky130_fd_sc_hd__xor2_1
XFILLER_178_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ rbzero.wall_tracer.visualWallDist\[-4\] _07252_ vssd1 vssd1 vccd1 vccd1 _07274_
+ sky130_fd_sc_hd__or2_1
XFILLER_53_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11829_ _03929_ _04540_ _04541_ _04542_ _03945_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__o221a_1
X_18385_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[3\] rbzero.spi_registers.spi_cmd\[2\]
+ rbzero.spi_registers.spi_cmd\[0\] vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__and4bb_1
X_15597_ _08193_ _08209_ _08210_ vssd1 vssd1 vccd1 vccd1 _08211_ sky130_fd_sc_hd__a21o_1
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17336_ _09744_ _09746_ vssd1 vssd1 vccd1 vccd1 _09875_ sky130_fd_sc_hd__nor2_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14548_ _07094_ _07219_ _07214_ _07085_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_187_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17267_ _09804_ _09805_ vssd1 vssd1 vccd1 vccd1 _09806_ sky130_fd_sc_hd__nor2_1
X_14479_ _07159_ _07061_ _07161_ _07163_ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__o22a_2
XFILLER_31_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19006_ rbzero.pov.spi_buffer\[50\] rbzero.pov.ready_buffer\[50\] _02662_ vssd1 vssd1
+ vccd1 vccd1 _02664_ sky130_fd_sc_hd__mux2_1
X_16218_ _08829_ _07410_ _07343_ vssd1 vssd1 vccd1 vccd1 _08830_ sky130_fd_sc_hd__mux2_1
X_17198_ _09606_ _09613_ _09612_ vssd1 vssd1 vccd1 vccd1 _09738_ sky130_fd_sc_hd__a21oi_1
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16149_ _07469_ _08760_ _08605_ _08602_ vssd1 vssd1 vccd1 vccd1 _08761_ sky130_fd_sc_hd__o31a_1
XFILLER_115_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19908_ _03113_ vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__clkinv_2
XFILLER_233_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19839_ _03107_ vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__clkinv_2
XFILLER_217_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20614_ net99 _00630_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20545_ net137 _00561_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20476_ net96 _00492_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21028_ net110 _01044_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13850_ _06317_ _06483_ vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__or2_1
XFILLER_142_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12801_ _05344_ _05357_ _05429_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__mux2_1
XFILLER_142_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13781_ _05660_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__buf_2
X_10993_ rbzero.tex_b0\[3\] rbzero.tex_b0\[2\] _03715_ vssd1 vssd1 vccd1 vccd1 _03725_
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15520_ _08084_ _08087_ vssd1 vssd1 vccd1 vccd1 _08134_ sky130_fd_sc_hd__xnor2_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _05361_ _05323_ _05325_ _05420_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__or4_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15451_ _07567_ _08060_ _08064_ _08063_ vssd1 vssd1 vccd1 vccd1 _08065_ sky130_fd_sc_hd__o31a_1
XFILLER_163_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _05341_ _05338_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__nor2_2
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14402_ _05401_ _06988_ _06985_ _05531_ vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__a211oi_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18170_ _01948_ _01949_ vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__or2b_1
XFILLER_187_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11614_ rbzero.tex_g0\[9\] rbzero.tex_g0\[8\] _04148_ vssd1 vssd1 vccd1 vccd1 _04331_
+ sky130_fd_sc_hd__mux2_1
X_15382_ _07995_ _07990_ vssd1 vssd1 vccd1 vccd1 _07996_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12594_ _03816_ _05069_ _05112_ _05282_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__a31o_1
XFILLER_145_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17121_ _09545_ _09561_ _09559_ vssd1 vssd1 vccd1 vccd1 _09661_ sky130_fd_sc_hd__a21o_1
XFILLER_168_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14333_ _07018_ _07021_ vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__or2b_1
XFILLER_141_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11545_ rbzero.debug_overlay.vplaneY\[-7\] _04238_ _04244_ rbzero.debug_overlay.vplaneY\[-1\]
+ _04246_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__a221o_1
XFILLER_106_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17052_ _08046_ _09055_ vssd1 vssd1 vccd1 vccd1 _09593_ sky130_fd_sc_hd__nand2_1
XFILLER_221_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14264_ _06927_ _06930_ _06908_ vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__a21oi_1
XFILLER_176_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11476_ _04192_ _04193_ _04099_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__mux2_1
XFILLER_143_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16003_ _08472_ _08480_ _08479_ vssd1 vssd1 vccd1 vccd1 _08616_ sky130_fd_sc_hd__a21bo_1
XFILLER_171_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13215_ _05883_ _05884_ _05902_ _05903_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__o31a_1
X_10427_ _03426_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__clkbuf_1
X_14195_ _06435_ _06634_ _06882_ _06883_ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__o31a_1
XFILLER_139_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13146_ _05827_ _05828_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__nand2_1
X_10358_ _03390_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17954_ _01588_ _01620_ _01628_ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__a21bo_2
X_13077_ _05635_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__inv_2
XFILLER_111_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10289_ _03353_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_239_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16905_ _09047_ _09188_ vssd1 vssd1 vccd1 vccd1 _09447_ sky130_fd_sc_hd__nor2_1
XFILLER_152_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12028_ _04735_ _04736_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__or2_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17885_ _01666_ _01667_ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__and2_1
XFILLER_22_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16836_ _09376_ _09377_ vssd1 vssd1 vccd1 vccd1 _09378_ sky130_fd_sc_hd__or2_1
X_19624_ _02834_ _02994_ _02995_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__or3_1
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19555_ _02946_ vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16767_ rbzero.wall_tracer.trackDistX\[-8\] _09301_ _09310_ _09316_ vssd1 vssd1 vccd1
+ vccd1 _00545_ sky130_fd_sc_hd__o22a_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13979_ _06101_ _06331_ _06320_ _06667_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18506_ _02191_ rbzero.debug_overlay.vplaneX\[-5\] vssd1 vssd1 vccd1 vccd1 _02252_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_207_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15718_ _08300_ _08303_ vssd1 vssd1 vccd1 vccd1 _08332_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19486_ rbzero.pov.spi_buffer\[39\] rbzero.pov.spi_buffer\[40\] _02910_ vssd1 vssd1
+ vccd1 vccd1 _02911_ sky130_fd_sc_hd__mux2_1
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16698_ rbzero.traced_texa\[0\] _09264_ _09265_ rbzero.wall_tracer.visualWallDist\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__a22o_1
XFILLER_179_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18437_ rbzero.debug_overlay.vplaneX\[-6\] _02170_ vssd1 vssd1 vccd1 vccd1 _02188_
+ sky130_fd_sc_hd__or2_1
X_15649_ _08237_ _08238_ vssd1 vssd1 vccd1 vccd1 _08263_ sky130_fd_sc_hd__xor2_1
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18368_ rbzero.wall_tracer.trackDistY\[9\] rbzero.wall_tracer.stepDistY\[9\] vssd1
+ vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__nand2_1
XFILLER_187_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17319_ _09728_ _09857_ vssd1 vssd1 vccd1 vccd1 _09858_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18299_ _02064_ _02065_ _02066_ _02061_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__o211a_1
XFILLER_30_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20330_ gpout1.clk_div\[0\] gpout1.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__or2_1
XFILLER_190_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20261_ _03125_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__buf_4
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20192_ _03211_ _03212_ _03213_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__a21o_1
XFILLER_66_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11330_ rbzero.row_render.size\[8\] rbzero.row_render.size\[7\] rbzero.row_render.size\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__nand3_1
XFILLER_193_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20528_ net120 _00544_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11261_ _03935_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__buf_4
X_20459_ net118 _00009_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13000_ _05607_ _05610_ _05619_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10212_ _03313_ vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11192_ _03905_ _03906_ _03910_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__mux2_1
XFILLER_238_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14951_ _07494_ _07564_ _07374_ vssd1 vssd1 vccd1 vccd1 _07565_ sky130_fd_sc_hd__mux2_1
XFILLER_48_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13902_ _06230_ _06176_ _06387_ _06529_ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__a31o_1
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17670_ _07886_ _10095_ _01454_ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__or3_1
XTAP_5887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14882_ rbzero.wall_tracer.visualWallDist\[0\] _03794_ vssd1 vssd1 vccd1 vccd1 _07496_
+ sky130_fd_sc_hd__nand2_1
XFILLER_235_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16621_ _09093_ _09091_ vssd1 vssd1 vccd1 vccd1 _09230_ sky130_fd_sc_hd__and2b_1
XFILLER_29_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13833_ _06440_ _06510_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__nor2_1
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19340_ _02857_ vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__clkinv_2
XFILLER_90_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16552_ _09024_ _09031_ _09160_ vssd1 vssd1 vccd1 vccd1 _09161_ sky130_fd_sc_hd__a21o_1
XFILLER_216_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13764_ _06450_ _06452_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__nand2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _03716_ vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15503_ _07416_ _07593_ vssd1 vssd1 vccd1 vccd1 _08117_ sky130_fd_sc_hd__nor2_1
X_12715_ _05360_ _05398_ _05401_ _05403_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__and4_2
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19271_ rbzero.spi_registers.new_other\[7\] rbzero.spi_registers.spi_buffer\[7\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__mux2_1
XFILLER_231_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16483_ _08846_ _08952_ _09092_ vssd1 vssd1 vccd1 vccd1 _09093_ sky130_fd_sc_hd__a21oi_1
XFILLER_188_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13695_ _06380_ _06382_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__nor2_1
XFILLER_245_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18222_ _02000_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__clkbuf_4
X_15434_ _07416_ _07508_ vssd1 vssd1 vccd1 vccd1 _08048_ sky130_fd_sc_hd__or2_1
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12646_ _05331_ _05332_ _05333_ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__or4_2
XFILLER_129_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18153_ _01730_ _01851_ _01731_ vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__o21ba_1
XFILLER_200_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15365_ _07975_ _07977_ vssd1 vssd1 vccd1 vccd1 _07979_ sky130_fd_sc_hd__or2b_1
X_12577_ _05175_ _05214_ _05174_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__a21bo_1
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17104_ _09642_ _09643_ _09644_ vssd1 vssd1 vccd1 vccd1 _09645_ sky130_fd_sc_hd__a21o_1
XFILLER_106_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14316_ _06987_ _06995_ _07004_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__o21ai_1
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18084_ _01863_ _01864_ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__xor2_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11528_ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__inv_2
X_15296_ _07517_ _07529_ _07620_ rbzero.wall_tracer.visualWallDist\[4\] vssd1 vssd1
+ vccd1 vccd1 _07910_ sky130_fd_sc_hd__or4b_1
XFILLER_183_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17035_ _07696_ _08640_ _07800_ vssd1 vssd1 vccd1 vccd1 _09576_ sky130_fd_sc_hd__a21o_1
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14247_ _06915_ _06917_ vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11459_ _04175_ _04176_ _03916_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__mux2_1
XFILLER_171_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14178_ _06865_ _06866_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__or2b_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13129_ _05706_ _05707_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__nand2_2
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _02653_ vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17937_ _01713_ _01718_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__nand2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17868_ _01567_ _01581_ _01650_ vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__a21bo_1
XFILLER_187_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19607_ rbzero.debug_overlay.playerX\[0\] _07562_ vssd1 vssd1 vccd1 vccd1 _02982_
+ sky130_fd_sc_hd__or2_1
XFILLER_113_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16819_ rbzero.wall_tracer.trackDistX\[-1\] rbzero.wall_tracer.stepDistX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _09362_ sky130_fd_sc_hd__nor2_1
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17799_ _01566_ _01582_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19538_ rbzero.pov.spi_buffer\[64\] rbzero.pov.spi_buffer\[65\] _02932_ vssd1 vssd1
+ vccd1 vccd1 _02938_ sky130_fd_sc_hd__mux2_1
XFILLER_59_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19469_ rbzero.pov.spi_buffer\[31\] rbzero.pov.spi_buffer\[32\] _02899_ vssd1 vssd1
+ vccd1 vccd1 _02902_ sky130_fd_sc_hd__mux2_1
XFILLER_107_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21362_ _00385_ _01378_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20313_ _08828_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__inv_2
XFILLER_200_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21293_ net134 _01309_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20244_ _03253_ vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__clkinv_2
XFILLER_235_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20175_ rbzero.traced_texa\[1\] rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1 _03200_
+ sky130_fd_sc_hd__nand2_1
XFILLER_27_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10830_ rbzero.tex_g0\[17\] rbzero.tex_g0\[16\] _03638_ vssd1 vssd1 vccd1 vccd1 _03640_
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10761_ rbzero.tex_g0\[49\] rbzero.tex_g0\[48\] _03593_ vssd1 vssd1 vccd1 vccd1 _03603_
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12500_ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__inv_2
XFILLER_197_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13480_ _06148_ _06150_ _06153_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__and3_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10692_ _03567_ vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12431_ _03733_ _05114_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__or2_1
XFILLER_201_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15150_ _07758_ _07763_ vssd1 vssd1 vccd1 vccd1 _07764_ sky130_fd_sc_hd__xor2_1
XFILLER_172_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12362_ _05053_ _05054_ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__and2_1
XFILLER_165_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14101_ _06632_ _06685_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__xor2_1
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11313_ _03902_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__buf_4
X_15081_ _07337_ _07688_ _07691_ _07694_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__o31a_2
X_12293_ _04959_ _04946_ _04986_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__nand3b_1
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14032_ _06669_ _06719_ vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__and2_1
XFILLER_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11244_ rbzero.tex_r0\[46\] _03962_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__and2_1
XFILLER_107_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11175_ _03893_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__buf_4
X_18840_ _02555_ _02556_ _02557_ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__o21a_1
XTAP_7075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18771_ _02468_ _02481_ _02482_ _02493_ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__o22a_1
XFILLER_95_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15983_ _08592_ vssd1 vssd1 vccd1 vccd1 _08596_ sky130_fd_sc_hd__buf_2
XTAP_5640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17722_ rbzero.wall_tracer.trackDistX\[6\] rbzero.wall_tracer.stepDistX\[6\] vssd1
+ vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__nor2_1
XTAP_5662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14934_ _07356_ _07547_ vssd1 vssd1 vccd1 vccd1 _07548_ sky130_fd_sc_hd__nand2_1
XFILLER_23_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17653_ _01430_ _01437_ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__xnor2_1
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14865_ _05093_ _05242_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__mux2_1
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16604_ _09211_ _09212_ vssd1 vssd1 vccd1 vccd1 _09213_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13816_ _06501_ _06499_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__xor2_1
X_17584_ _09861_ _09989_ _10120_ vssd1 vssd1 vccd1 vccd1 _10121_ sky130_fd_sc_hd__o21a_2
XFILLER_223_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14796_ rbzero.debug_overlay.playerX\[-4\] vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__inv_2
XFILLER_56_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19323_ _02852_ _02853_ vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__nor2_1
X_16535_ _08086_ _07597_ _07621_ _08223_ vssd1 vssd1 vccd1 vccd1 _09144_ sky130_fd_sc_hd__o22a_1
XFILLER_232_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13747_ _06376_ _06379_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__and2_1
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10959_ _03707_ vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19254_ _02810_ vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16466_ _09071_ _09072_ _09074_ vssd1 vssd1 vccd1 vccd1 _09076_ sky130_fd_sc_hd__a21o_1
XFILLER_231_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13678_ _06323_ _06364_ _06366_ vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__o21a_1
X_18205_ _01981_ _01984_ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__xnor2_1
X_15417_ _08027_ _08029_ _08030_ vssd1 vssd1 vccd1 vccd1 _08031_ sky130_fd_sc_hd__a21oi_1
XFILLER_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12629_ _05315_ _05317_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__xor2_1
X_19185_ rbzero.spi_registers.new_floor\[4\] rbzero.color_floor\[4\] _02763_ vssd1
+ vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__mux2_1
X_16397_ _09003_ _09005_ vssd1 vssd1 vccd1 vccd1 _09007_ sky130_fd_sc_hd__and2_1
XFILLER_157_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18136_ _01824_ _01826_ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__nand2_1
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15348_ _07613_ _07612_ vssd1 vssd1 vccd1 vccd1 _07962_ sky130_fd_sc_hd__and2b_1
XFILLER_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18067_ _01736_ _01847_ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15279_ _07424_ _07567_ vssd1 vssd1 vccd1 vccd1 _07893_ sky130_fd_sc_hd__or2_1
XFILLER_144_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17018_ _09556_ _09558_ vssd1 vssd1 vccd1 vccd1 _09559_ sky130_fd_sc_hd__nor2_1
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18969_ _02644_ vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20931_ net74 _00947_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[68\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20862_ _00080_ _00878_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[63\] sky130_fd_sc_hd__dfxtp_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20793_ net86 _00809_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21345_ _00368_ _01361_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21276_ _00325_ _01292_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20227_ _03240_ _03241_ _03242_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__nand3_1
XFILLER_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20158_ _03184_ _03185_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__xor2_1
XFILLER_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12980_ _05624_ _05660_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__nor2_1
X_20089_ _03131_ vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__clkinv_2
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11931_ _04615_ _04638_ _04640_ _04641_ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__and4_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14650_ rbzero.wall_tracer.visualWallDist\[6\] _07252_ vssd1 vssd1 vccd1 vccd1 _07297_
+ sky130_fd_sc_hd__or2_1
XFILLER_150_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _03909_ _04573_ _04574_ _04575_ _03944_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__o221a_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _06224_ _06258_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__and2_1
XFILLER_150_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10813_ rbzero.tex_g0\[25\] rbzero.tex_g0\[24\] _03627_ vssd1 vssd1 vccd1 vccd1 _03631_
+ sky130_fd_sc_hd__mux2_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14581_ _05025_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__clkbuf_4
XFILLER_26_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11793_ _04506_ _04507_ _03916_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__mux2_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16320_ _08929_ _08930_ vssd1 vssd1 vccd1 vccd1 _08931_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13532_ _06218_ _06220_ vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__xor2_1
XFILLER_207_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10744_ _03594_ vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16251_ _08853_ _08861_ vssd1 vssd1 vccd1 vccd1 _08862_ sky130_fd_sc_hd__xnor2_1
XFILLER_186_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13463_ _05981_ _06022_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10675_ _03558_ vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15202_ _07455_ _07641_ vssd1 vssd1 vccd1 vccd1 _07816_ sky130_fd_sc_hd__and2_1
XFILLER_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12414_ _05064_ _05057_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__nor2_1
X_16182_ _07824_ _08793_ _07835_ vssd1 vssd1 vccd1 vccd1 _08794_ sky130_fd_sc_hd__a21o_1
XFILLER_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13394_ _06071_ _06073_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__nand2_1
XFILLER_194_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15133_ _07727_ _07737_ _07725_ vssd1 vssd1 vccd1 vccd1 _07747_ sky130_fd_sc_hd__a21bo_1
XFILLER_126_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12345_ rbzero.debug_overlay.facingY\[-7\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__or2_1
XFILLER_177_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15064_ _04929_ _07651_ vssd1 vssd1 vccd1 vccd1 _07678_ sky130_fd_sc_hd__nand2_1
XFILLER_173_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19941_ _03117_ vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__clkinv_2
X_12276_ _04968_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.trackDistY\[-12\]
+ _04969_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__o22a_1
XFILLER_181_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14015_ _06636_ _06638_ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__or2_1
X_11227_ _03945_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__clkbuf_4
X_19872_ _03110_ vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__clkinv_2
XFILLER_229_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18823_ _03819_ _02532_ _02533_ _02542_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__a31o_1
XTAP_6160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11158_ rbzero.texV\[7\] _03832_ _03830_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__a21oi_1
XTAP_6171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15966_ _08573_ _08575_ vssd1 vssd1 vccd1 vccd1 _08580_ sky130_fd_sc_hd__nor2_1
X_18754_ _02475_ _02476_ _02473_ _02474_ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__o211ai_2
X_11089_ _03811_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__clkbuf_4
XFILLER_209_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17705_ _10090_ _10132_ _01489_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__a21oi_1
XFILLER_188_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14917_ _07524_ _07529_ _07523_ vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15897_ _07598_ _08510_ vssd1 vssd1 vccd1 vccd1 _08511_ sky130_fd_sc_hd__nor2_1
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18685_ rbzero.debug_overlay.vplaneY\[-6\] _02396_ vssd1 vssd1 vccd1 vccd1 _02414_
+ sky130_fd_sc_hd__or2_1
XFILLER_236_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17636_ _09166_ _08723_ vssd1 vssd1 vccd1 vccd1 _10172_ sky130_fd_sc_hd__or2_1
X_14848_ rbzero.debug_overlay.playerX\[-7\] vssd1 vssd1 vccd1 vccd1 _07462_ sky130_fd_sc_hd__inv_2
XFILLER_64_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17567_ _09836_ _09961_ vssd1 vssd1 vccd1 vccd1 _10104_ sky130_fd_sc_hd__nand2_1
XFILLER_225_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14779_ rbzero.wall_tracer.visualWallDist\[-5\] _03793_ vssd1 vssd1 vccd1 vccd1 _07393_
+ sky130_fd_sc_hd__and2_1
XFILLER_229_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16518_ _08429_ _08979_ vssd1 vssd1 vccd1 vccd1 _09127_ sky130_fd_sc_hd__nor2_1
X_19306_ rbzero.pov.spi_counter\[0\] _02837_ rbzero.pov.spi_counter\[1\] vssd1 vssd1
+ vccd1 vccd1 _02841_ sky130_fd_sc_hd__a21o_1
XFILLER_232_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17498_ _10018_ vssd1 vssd1 vccd1 vccd1 _10035_ sky130_fd_sc_hd__inv_2
XFILLER_225_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16449_ _09056_ _09057_ _09058_ vssd1 vssd1 vccd1 vccd1 _09059_ sky130_fd_sc_hd__nand3_1
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19237_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.new_floor\[5\]
+ _02795_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__mux2_1
XFILLER_176_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19168_ _02759_ vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__clkbuf_1
XFILLER_157_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18119_ _01805_ _01899_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19099_ _02713_ vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21130_ _00179_ _01146_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21061_ _00110_ _01077_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20012_ _03123_ vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__clkinv_2
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20914_ net74 _00930_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[51\] sky130_fd_sc_hd__dfxtp_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20845_ _00063_ _00861_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_243_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20776_ net88 _00792_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout55 net57 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_2
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout66 net72 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_2
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout77 net78 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout88 net89 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout99 net100 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_2
XFILLER_211_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10460_ _03444_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__clkbuf_4
XFILLER_52_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10391_ _03407_ vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12130_ _03288_ gpout0.hpos\[1\] _04631_ _04632_ net27 _04832_ vssd1 vssd1 vccd1
+ vccd1 _04837_ sky130_fd_sc_hd__mux4_1
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21328_ _00351_ _01344_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12061_ _04768_ _04447_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__nand2_1
X_21259_ _00308_ _01275_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11012_ _03736_ _03733_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__xor2_1
XFILLER_78_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15820_ _08428_ _08398_ _08426_ _08433_ vssd1 vssd1 vccd1 vccd1 _08434_ sky130_fd_sc_hd__or4bb_1
XFILLER_172_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _07880_ _08336_ _08136_ _08337_ vssd1 vssd1 vccd1 vccd1 _08365_ sky130_fd_sc_hd__and4bb_1
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12963_ _05624_ _05622_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__nor2_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _07325_ vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__clkbuf_1
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11914_ net14 net13 _04624_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__and3_1
X_18470_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__nand2_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15682_ _08295_ vssd1 vssd1 vccd1 vccd1 _08296_ sky130_fd_sc_hd__buf_4
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12894_ _05582_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__inv_2
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _07886_ _09829_ vssd1 vssd1 vccd1 vccd1 _09959_ sky130_fd_sc_hd__nor2_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ rbzero.wall_tracer.visualWallDist\[1\] _07252_ vssd1 vssd1 vccd1 vccd1 _07285_
+ sky130_fd_sc_hd__or2_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11845_ _04557_ _04558_ _03908_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__mux2_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _09766_ _09770_ vssd1 vssd1 vccd1 vccd1 _09891_ sky130_fd_sc_hd__nand2_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14564_ _05408_ _07231_ _07232_ _07075_ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__o211a_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ rbzero.tex_b0\[17\] rbzero.tex_b0\[16\] _04001_ vssd1 vssd1 vccd1 vccd1 _04491_
+ sky130_fd_sc_hd__mux2_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _08912_ _08913_ vssd1 vssd1 vccd1 vccd1 _08914_ sky130_fd_sc_hd__nor2_1
XFILLER_207_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13515_ _06196_ _06197_ _06203_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__o21ai_1
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17283_ _09820_ _09821_ vssd1 vssd1 vccd1 vccd1 _09822_ sky130_fd_sc_hd__nor2_1
XFILLER_186_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10727_ _03585_ vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14495_ _07107_ _07139_ _07177_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__a21o_1
X_19022_ rbzero.pov.spi_buffer\[58\] rbzero.pov.ready_buffer\[58\] _02662_ vssd1 vssd1
+ vccd1 vccd1 _02672_ sky130_fd_sc_hd__mux2_1
X_16234_ _08841_ _08843_ vssd1 vssd1 vccd1 vccd1 _08845_ sky130_fd_sc_hd__and2_1
XFILLER_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13446_ _06126_ _06134_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__nand2_1
X_10658_ _03549_ vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16165_ _08770_ _08776_ vssd1 vssd1 vccd1 vccd1 _08777_ sky130_fd_sc_hd__xnor2_1
XFILLER_103_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13377_ _06061_ _06062_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__xor2_1
X_10589_ _03513_ vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15116_ _07213_ _07195_ _07346_ vssd1 vssd1 vccd1 vccd1 _07730_ sky130_fd_sc_hd__a21o_1
XFILLER_155_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12328_ _05019_ _04989_ _05021_ _04967_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__or4b_1
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16096_ rbzero.wall_tracer.texu\[1\] _07338_ _08707_ _08708_ _07266_ vssd1 vssd1
+ vccd1 vccd1 _00482_ sky130_fd_sc_hd__o221a_1
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15047_ _04932_ _07658_ _07660_ _07453_ vssd1 vssd1 vccd1 vccd1 _07661_ sky130_fd_sc_hd__a211o_1
XFILLER_170_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19924_ _03115_ vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__clkinv_2
X_12259_ rbzero.wall_tracer.trackDistY\[-1\] vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__inv_2
XFILLER_218_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19855_ _03108_ vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__clkinv_2
XFILLER_151_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18806_ rbzero.wall_tracer.rayAddendY\[6\] _02197_ _02526_ _02166_ vssd1 vssd1 vccd1
+ vccd1 _02527_ sky130_fd_sc_hd__a22o_1
X_19786_ _03090_ vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16998_ _08599_ _08724_ vssd1 vssd1 vccd1 vccd1 _09539_ sky130_fd_sc_hd__nor2_1
XFILLER_209_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18737_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.debug_overlay.vplaneY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__nor2_1
XFILLER_237_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15949_ _08561_ _08562_ vssd1 vssd1 vccd1 vccd1 _08563_ sky130_fd_sc_hd__and2_2
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18668_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.wall_tracer.rayAddendY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__nor2_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17619_ _10065_ _10068_ _10154_ vssd1 vssd1 vccd1 vccd1 _10155_ sky130_fd_sc_hd__a21o_1
XFILLER_224_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18599_ _02327_ _02330_ _02337_ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20630_ net56 _00646_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20561_ net136 _00577_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20492_ net114 _00508_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21113_ _00162_ _01129_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_6907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21044_ _00093_ _01060_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ rbzero.tex_g0\[57\] rbzero.tex_g0\[56\] _04000_ vssd1 vssd1 vccd1 vccd1 _04347_
+ sky130_fd_sc_hd__mux2_1
X_20828_ _00046_ _00844_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11561_ rbzero.debug_overlay.playerY\[3\] _04231_ _04244_ rbzero.debug_overlay.playerY\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__a22o_1
XFILLER_243_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20759_ net107 _00775_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13300_ _05984_ _05988_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__and2_1
XFILLER_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10512_ rbzero.tex_r0\[40\] rbzero.tex_r0\[39\] _03468_ vssd1 vssd1 vccd1 vccd1 _03473_
+ sky130_fd_sc_hd__mux2_1
X_14280_ _06791_ _06967_ _06968_ vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__o21ba_1
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11492_ gpout0.hpos\[5\] _03806_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__xor2_1
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13231_ _05918_ _05889_ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__nor3_1
XFILLER_100_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10443_ rbzero.tex_r1\[6\] rbzero.tex_r1\[7\] _03433_ vssd1 vssd1 vccd1 vccd1 _03435_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13162_ _05849_ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__or2_1
XFILLER_164_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10374_ _03398_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12113_ net27 vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__buf_2
XFILLER_112_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17970_ _01736_ _01751_ vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__xnor2_1
X_13093_ _05721_ _05733_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__nand2_1
XFILLER_124_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16921_ _09462_ vssd1 vssd1 vccd1 vccd1 _09463_ sky130_fd_sc_hd__clkbuf_4
X_12044_ net7 net8 vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__and2b_1
XFILLER_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19640_ rbzero.debug_overlay.playerY\[-9\] vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__inv_2
XFILLER_120_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16852_ _09392_ _09393_ vssd1 vssd1 vccd1 vccd1 _09394_ sky130_fd_sc_hd__nand2_1
XFILLER_238_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15803_ _08356_ _08382_ vssd1 vssd1 vccd1 vccd1 _08417_ sky130_fd_sc_hd__and2_1
XFILLER_133_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16783_ rbzero.wall_tracer.trackDistX\[-6\] _09301_ _09324_ _09330_ vssd1 vssd1 vccd1
+ vccd1 _00547_ sky130_fd_sc_hd__o22a_1
X_19571_ net39 _02954_ _02721_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__o21ai_4
XFILLER_24_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13995_ _06681_ _06683_ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__or2b_1
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15734_ _08331_ _08347_ vssd1 vssd1 vccd1 vccd1 _08348_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18522_ _02266_ _02252_ _02238_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__a21bo_1
X_12946_ _05545_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__clkbuf_4
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15665_ _08232_ _08236_ vssd1 vssd1 vccd1 vccd1 _08279_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18453_ _09261_ _02195_ _02196_ _02202_ vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__a31o_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12877_ _05526_ _05546_ _05553_ _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__a31o_1
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17404_ _09808_ _09817_ _09815_ vssd1 vssd1 vccd1 vccd1 _09942_ sky130_fd_sc_hd__a21oi_1
X_14616_ rbzero.wall_tracer.trackDistX\[-4\] rbzero.wall_tracer.trackDistY\[-4\] _07258_
+ vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__mux2_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18384_ _01990_ _02139_ _01996_ rbzero.wall_tracer.trackDistY\[11\] vssd1 vssd1 vccd1
+ vccd1 _00588_ sky130_fd_sc_hd__o2bb2a_1
X_11828_ rbzero.tex_b1\[41\] _03938_ _03940_ _03908_ vssd1 vssd1 vccd1 vccd1 _04542_
+ sky130_fd_sc_hd__a31o_1
X_15596_ _08194_ _08208_ vssd1 vssd1 vccd1 vccd1 _08210_ sky130_fd_sc_hd__nor2_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17335_ _09825_ _09873_ vssd1 vssd1 vccd1 vccd1 _09874_ sky130_fd_sc_hd__xnor2_1
XFILLER_226_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _05568_ _07007_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__nor2_1
XFILLER_187_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11759_ _04472_ _04473_ _03916_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__mux2_1
XFILLER_159_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17266_ _09802_ _09803_ vssd1 vssd1 vccd1 vccd1 _09805_ sky130_fd_sc_hd__and2_1
XFILLER_201_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14478_ _05447_ _07162_ _05602_ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__a21o_1
XFILLER_140_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16217_ rbzero.debug_overlay.playerY\[-4\] vssd1 vssd1 vccd1 vccd1 _08829_ sky130_fd_sc_hd__clkinv_2
X_19005_ _02663_ vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13429_ _06116_ _06117_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__xnor2_1
X_17197_ _09730_ _09736_ vssd1 vssd1 vccd1 vccd1 _09737_ sky130_fd_sc_hd__xor2_1
XFILLER_220_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16148_ _07805_ vssd1 vssd1 vccd1 vccd1 _08760_ sky130_fd_sc_hd__clkbuf_4
XFILLER_31_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16079_ _07628_ _07921_ _08550_ _08548_ vssd1 vssd1 vccd1 vccd1 _08692_ sky130_fd_sc_hd__o31a_1
XFILLER_130_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19907_ _03113_ vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__clkinv_2
XFILLER_216_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19838_ _03107_ vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__clkinv_2
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput1 i_clk vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_6
X_19769_ o_vsync _03075_ _03077_ vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__a21boi_1
XFILLER_232_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20613_ net99 _00629_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_240_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20544_ net137 _00560_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20475_ net96 _00491_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_119_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21027_ net109 _01043_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12800_ _05471_ _05474_ _05488_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__a21o_2
X_13780_ _05651_ _06311_ _06468_ _05434_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__a211o_1
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10992_ _03724_ vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12731_ _05327_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__inv_2
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ _08061_ _08062_ _08063_ vssd1 vssd1 vccd1 vccd1 _08064_ sky130_fd_sc_hd__a21bo_1
XFILLER_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12662_ _05323_ _05325_ _05327_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__or3_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14401_ _07075_ _07086_ _07089_ vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__or3b_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _04328_ _04329_ _04014_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__mux2_1
XFILLER_93_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15381_ _07610_ _07983_ vssd1 vssd1 vccd1 vccd1 _07995_ sky130_fd_sc_hd__nor2_1
XFILLER_212_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12593_ rbzero.wall_tracer.visualWallDist\[4\] _05190_ vssd1 vssd1 vccd1 vccd1 _05282_
+ sky130_fd_sc_hd__and2_1
XFILLER_204_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17120_ _09520_ _09659_ vssd1 vssd1 vccd1 vccd1 _09660_ sky130_fd_sc_hd__xor2_1
XFILLER_141_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14332_ _06981_ _07020_ vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__nand2_1
XFILLER_180_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11544_ rbzero.debug_overlay.vplaneY\[-3\] _04209_ _04243_ rbzero.debug_overlay.vplaneY\[0\]
+ _04261_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__a221o_1
XFILLER_102_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17051_ _09449_ _09197_ _09188_ vssd1 vssd1 vccd1 vccd1 _09592_ sky130_fd_sc_hd__or3_1
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14263_ _06931_ _06944_ _06950_ _06951_ vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__and4_1
XFILLER_184_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11475_ rbzero.color_sky\[1\] rbzero.color_floor\[1\] _04030_ vssd1 vssd1 vccd1 vccd1
+ _04193_ sky130_fd_sc_hd__mux2_1
XFILLER_221_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16002_ _07858_ _07736_ _08465_ _08464_ vssd1 vssd1 vccd1 vccd1 _08615_ sky130_fd_sc_hd__o31ai_1
XFILLER_137_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13214_ _05901_ _05885_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__or2b_1
X_10426_ rbzero.tex_r1\[14\] rbzero.tex_r1\[15\] _03422_ vssd1 vssd1 vccd1 vccd1 _03426_
+ sky130_fd_sc_hd__mux2_1
X_14194_ _06137_ _06343_ _06881_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__or3_1
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13145_ _05832_ _05833_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10357_ rbzero.tex_r1\[47\] rbzero.tex_r1\[48\] _03389_ vssd1 vssd1 vccd1 vccd1 _03390_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _01635_ _01642_ _01734_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__a21o_1
X_13076_ _05763_ _05764_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__or2_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10288_ rbzero.tex_b1\[15\] rbzero.tex_b1\[16\] _03344_ vssd1 vssd1 vccd1 vccd1 _03353_
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16904_ _09425_ _09445_ vssd1 vssd1 vccd1 vccd1 _09446_ sky130_fd_sc_hd__xnor2_1
X_12027_ _03288_ gpout0.hpos\[1\] gpout0.vpos\[0\] _04632_ net3 _04731_ vssd1 vssd1
+ vccd1 vccd1 _04736_ sky130_fd_sc_hd__mux4_1
XFILLER_215_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17884_ _01656_ _01665_ vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__or2_1
XFILLER_152_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19623_ rbzero.debug_overlay.playerX\[3\] _02991_ vssd1 vssd1 vccd1 vccd1 _02995_
+ sky130_fd_sc_hd__nor2_1
XFILLER_113_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16835_ _09135_ _09138_ _09375_ vssd1 vssd1 vccd1 vccd1 _09377_ sky130_fd_sc_hd__and3_1
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19554_ rbzero.pov.spi_buffer\[72\] rbzero.pov.spi_buffer\[73\] _02865_ vssd1 vssd1
+ vccd1 vccd1 _02946_ sky130_fd_sc_hd__mux2_1
XFILLER_207_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13978_ _06470_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__clkinv_2
X_16766_ _09303_ _09314_ _09315_ _09283_ vssd1 vssd1 vccd1 vccd1 _09316_ sky130_fd_sc_hd__a31o_1
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18505_ _02248_ _02249_ _02245_ _02246_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__a211o_1
X_15717_ _08290_ _08306_ vssd1 vssd1 vccd1 vccd1 _08331_ sky130_fd_sc_hd__xnor2_1
X_12929_ _05617_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__buf_2
XFILLER_146_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16697_ _09257_ vssd1 vssd1 vccd1 vccd1 _09265_ sky130_fd_sc_hd__buf_2
X_19485_ _02865_ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__clkbuf_4
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18436_ rbzero.debug_overlay.vplaneX\[-6\] _02170_ vssd1 vssd1 vccd1 vccd1 _02187_
+ sky130_fd_sc_hd__nand2_1
X_15648_ _08251_ _08260_ _08261_ vssd1 vssd1 vccd1 vccd1 _08262_ sky130_fd_sc_hd__a21o_1
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18367_ rbzero.wall_tracer.trackDistY\[9\] rbzero.wall_tracer.stepDistY\[9\] vssd1
+ vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__or2_1
X_15579_ _08183_ _08184_ vssd1 vssd1 vccd1 vccd1 _08193_ sky130_fd_sc_hd__xor2_1
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17318_ _09465_ _09466_ _09732_ vssd1 vssd1 vccd1 vccd1 _09857_ sky130_fd_sc_hd__and3_1
XFILLER_174_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18298_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.stepDistY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__nand2_1
XFILLER_120_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17249_ _09656_ _09787_ vssd1 vssd1 vccd1 vccd1 _09788_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20260_ _03254_ vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__clkinv_2
XFILLER_200_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20191_ _03211_ _03212_ _03213_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__nand3_1
XFILLER_131_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20527_ net120 _00543_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11260_ rbzero.tex_r0\[35\] _03939_ _03941_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__and3_1
XFILLER_197_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20458_ net118 _00008_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10211_ rbzero.tex_b1\[52\] rbzero.tex_b1\[53\] _03311_ vssd1 vssd1 vccd1 vccd1 _03313_
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11191_ _03909_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__buf_4
XFILLER_79_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20389_ net135 _00420_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14950_ _07562_ _07563_ vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__nand2_1
XFILLER_212_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13901_ _06587_ _06588_ _06589_ vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__a21o_1
XFILLER_130_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14881_ _07492_ _07493_ _07494_ vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__and3b_1
XFILLER_43_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16620_ _08972_ _09228_ vssd1 vssd1 vccd1 vccd1 _09229_ sky130_fd_sc_hd__xnor2_1
X_13832_ _06519_ _06520_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__or2b_1
XFILLER_78_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16551_ _09029_ _09030_ vssd1 vssd1 vccd1 vccd1 _09160_ sky130_fd_sc_hd__nor2_1
XFILLER_204_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13763_ _06400_ _06451_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__and2_1
XFILLER_245_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10975_ rbzero.tex_b0\[12\] rbzero.tex_b0\[11\] _03715_ vssd1 vssd1 vccd1 vccd1 _03716_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12714_ _05328_ _05335_ _05402_ _05383_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__o211ai_1
X_15502_ _08093_ _08094_ vssd1 vssd1 vccd1 vccd1 _08116_ sky130_fd_sc_hd__xnor2_2
X_16482_ _08949_ _08951_ vssd1 vssd1 vccd1 vccd1 _09092_ sky130_fd_sc_hd__nor2_1
X_19270_ _02819_ vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__clkbuf_1
XFILLER_245_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13694_ _06380_ _06382_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__and2_1
XFILLER_206_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18221_ _03797_ _08629_ _05027_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__o21ai_2
XFILLER_176_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15433_ _08046_ _07579_ vssd1 vssd1 vccd1 vccd1 _08047_ sky130_fd_sc_hd__nand2_1
XFILLER_231_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12645_ _05296_ _05265_ _05270_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18152_ _01736_ _01931_ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__xnor2_1
X_15364_ _07975_ _07977_ vssd1 vssd1 vccd1 vccd1 _07978_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12576_ _05211_ _05213_ _05218_ _05224_ _05264_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a2111o_1
XFILLER_106_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14315_ _06985_ _07003_ vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__or2_1
X_17103_ rbzero.wall_tracer.trackDistX\[0\] rbzero.wall_tracer.stepDistX\[0\] _09511_
+ vssd1 vssd1 vccd1 vccd1 _09644_ sky130_fd_sc_hd__a21o_1
XFILLER_15_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18083_ _09829_ _08725_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__nor2_1
XFILLER_157_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11527_ gpout0.hpos\[4\] _04215_ _04233_ _03780_ vssd1 vssd1 vccd1 vccd1 _04245_
+ sky130_fd_sc_hd__and4bb_2
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15295_ _07811_ _07784_ vssd1 vssd1 vccd1 vccd1 _07909_ sky130_fd_sc_hd__or2b_1
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17034_ _09573_ _09574_ vssd1 vssd1 vccd1 vccd1 _09575_ sky130_fd_sc_hd__xnor2_2
XFILLER_32_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14246_ _06914_ _06934_ vssd1 vssd1 vccd1 vccd1 _06935_ sky130_fd_sc_hd__or2_1
XFILLER_172_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11458_ rbzero.tex_r1\[13\] rbzero.tex_r1\[12\] _04168_ vssd1 vssd1 vccd1 vccd1 _04176_
+ sky130_fd_sc_hd__mux2_1
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10409_ rbzero.tex_r1\[22\] rbzero.tex_r1\[23\] _03411_ vssd1 vssd1 vccd1 vccd1 _03417_
+ sky130_fd_sc_hd__mux2_1
X_14177_ _06857_ _06863_ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__xor2_1
XFILLER_139_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11389_ gpout0.vpos\[2\] gpout0.vpos\[1\] gpout0.vpos\[0\] _04107_ vssd1 vssd1 vccd1
+ vccd1 _04108_ sky130_fd_sc_hd__o31a_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13128_ _05815_ _05816_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__xor2_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ rbzero.pov.spi_buffer\[40\] rbzero.pov.ready_buffer\[40\] _02651_ vssd1 vssd1
+ vccd1 vccd1 _02653_ sky130_fd_sc_hd__mux2_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17936_ _01713_ _01718_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__nor2_1
X_13059_ _05564_ _05613_ _05614_ _05616_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__or4_4
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17867_ _01582_ _01566_ vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__or2b_1
XFILLER_22_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19606_ net39 _02954_ _02720_ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__o21a_1
X_16818_ _09351_ _09237_ vssd1 vssd1 vccd1 vccd1 _09361_ sky130_fd_sc_hd__nand2_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17798_ _01567_ _01581_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19537_ _02937_ vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__clkbuf_1
X_16749_ rbzero.wall_tracer.trackDistX\[-10\] _09276_ _09294_ _09300_ vssd1 vssd1
+ vccd1 vccd1 _00543_ sky130_fd_sc_hd__o22a_1
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19468_ _02901_ vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18419_ rbzero.debug_overlay.vplaneX\[-7\] _02168_ vssd1 vssd1 vccd1 vccd1 _02171_
+ sky130_fd_sc_hd__nand2_1
XFILLER_222_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19399_ _02838_ _02837_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__nand2_2
XFILLER_210_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21361_ _00384_ _01377_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20312_ _08700_ _09269_ rbzero.traced_texVinit\[3\] _09255_ vssd1 vssd1 vccd1 vccd1
+ _01397_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_194_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21292_ net134 _01308_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20243_ _03253_ vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__clkinv_2
XFILLER_107_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20174_ rbzero.traced_texa\[1\] rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1 _03199_
+ sky130_fd_sc_hd__or2_1
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10760_ _03602_ vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10691_ rbzero.tex_g1\[18\] rbzero.tex_g1\[19\] _03563_ vssd1 vssd1 vccd1 vccd1 _03567_
+ sky130_fd_sc_hd__mux2_1
XFILLER_205_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12430_ _03733_ _05114_ vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__nand2_1
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12361_ rbzero.debug_overlay.facingY\[-1\] rbzero.wall_tracer.rayAddendY\[7\] vssd1
+ vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__or2_1
XFILLER_51_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14100_ _06782_ _06788_ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__and2_1
XFILLER_193_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11312_ rbzero.color_sky\[0\] rbzero.color_floor\[0\] _04030_ vssd1 vssd1 vccd1 vccd1
+ _04031_ sky130_fd_sc_hd__mux2_1
X_15080_ _03794_ _07693_ vssd1 vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__and2_4
XFILLER_180_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12292_ _04985_ rbzero.wall_tracer.trackDistY\[3\] rbzero.wall_tracer.trackDistY\[-4\]
+ _04948_ _04943_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__o221a_1
XFILLER_153_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14031_ _06669_ _06719_ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__xor2_1
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11243_ _03961_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__clkbuf_4
XTAP_7021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11174_ _03891_ _03892_ rbzero.row_render.vinf vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__a21oi_1
XTAP_7076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18770_ _04260_ rbzero.debug_overlay.vplaneY\[-6\] vssd1 vssd1 vccd1 vccd1 _02493_
+ sky130_fd_sc_hd__nor2_1
XTAP_6375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15982_ _07790_ vssd1 vssd1 vccd1 vccd1 _08595_ sky130_fd_sc_hd__clkbuf_4
XTAP_5630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17721_ _01500_ _01503_ _01505_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__a21oi_2
XTAP_5663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14933_ _07493_ _07546_ _07374_ vssd1 vssd1 vccd1 vccd1 _07547_ sky130_fd_sc_hd__mux2_1
XTAP_5674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17652_ _01431_ _01436_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__xor2_1
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14864_ _07100_ _07171_ _07336_ vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__a21o_1
XFILLER_35_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16603_ _09056_ _09059_ vssd1 vssd1 vccd1 vccd1 _09212_ sky130_fd_sc_hd__nand2_1
X_13815_ _06456_ _06503_ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__xor2_1
XFILLER_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17583_ _09861_ _09988_ vssd1 vssd1 vccd1 vccd1 _10120_ sky130_fd_sc_hd__nand2_1
X_14795_ rbzero.wall_tracer.visualWallDist\[-4\] _07407_ _07408_ vssd1 vssd1 vccd1
+ vccd1 _07409_ sky130_fd_sc_hd__mux2_1
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19322_ rbzero.pov.spi_counter\[5\] _02849_ _02838_ vssd1 vssd1 vccd1 vccd1 _02853_
+ sky130_fd_sc_hd__o21ai_1
X_16534_ _08890_ _08671_ vssd1 vssd1 vccd1 vccd1 _09143_ sky130_fd_sc_hd__nor2_1
X_13746_ _05638_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__clkbuf_4
XFILLER_1_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10958_ rbzero.tex_b0\[20\] rbzero.tex_b0\[19\] _03704_ vssd1 vssd1 vccd1 vccd1 _03707_
+ sky130_fd_sc_hd__mux2_1
XFILLER_231_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19253_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.new_leak\[5\] _02804_
+ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__mux2_1
X_16465_ _09071_ _09072_ _09074_ vssd1 vssd1 vccd1 vccd1 _09075_ sky130_fd_sc_hd__nand3_1
XFILLER_188_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13677_ _06308_ _06365_ _06319_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__o21ai_1
XFILLER_189_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10889_ _03670_ vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18204_ _01896_ _01983_ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__xnor2_1
XPHY_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15416_ _08004_ _08026_ vssd1 vssd1 vccd1 vccd1 _08030_ sky130_fd_sc_hd__nor2_1
X_12628_ _05305_ _05312_ _05316_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__a21o_1
X_16396_ _09003_ _09005_ vssd1 vssd1 vccd1 vccd1 _09006_ sky130_fd_sc_hd__nor2_1
XFILLER_157_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19184_ rbzero.color_floor\[3\] _02763_ _02769_ vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__a21o_1
XPHY_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18135_ _05121_ _01914_ _01915_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__or3_2
X_15347_ _07640_ _07960_ vssd1 vssd1 vccd1 vccd1 _07961_ sky130_fd_sc_hd__xnor2_2
X_12559_ rbzero.wall_tracer.visualWallDist\[-8\] _05095_ rbzero.wall_tracer.rcp_sel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__mux2_1
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18066_ _01842_ _01846_ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__xnor2_1
X_15278_ _07889_ _07891_ vssd1 vssd1 vccd1 vccd1 _07892_ sky130_fd_sc_hd__nand2_1
XFILLER_176_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17017_ _09404_ _09412_ _09557_ vssd1 vssd1 vccd1 vccd1 _09558_ sky130_fd_sc_hd__a21oi_1
X_14229_ _06889_ _06914_ _06915_ _06917_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_217_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18968_ rbzero.pov.spi_buffer\[32\] rbzero.pov.ready_buffer\[32\] _02640_ vssd1 vssd1
+ vccd1 vccd1 _02644_ sky130_fd_sc_hd__mux2_1
XFILLER_227_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17919_ _01690_ _01701_ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__xnor2_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18899_ _02606_ vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__clkbuf_4
XFILLER_239_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20930_ net74 _00946_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[67\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20861_ _00079_ _00877_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20792_ net84 _00808_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_241_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21344_ _00367_ _01360_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21275_ _00324_ _01291_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20226_ _03240_ _03241_ _03242_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__a21o_1
XFILLER_46_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20157_ _03177_ _03179_ _03178_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__a21boi_1
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20088_ _03131_ vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__clkinv_2
XFILLER_217_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11930_ net12 net13 _04639_ net14 vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__o22a_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11861_ rbzero.tex_b1\[10\] _03903_ _03928_ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a21o_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _06261_ _06288_ vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__xnor2_4
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10812_ _03630_ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _03799_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__buf_2
XFILLER_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11792_ rbzero.tex_b0\[13\] rbzero.tex_b0\[12\] _03925_ vssd1 vssd1 vccd1 vccd1 _04507_
+ sky130_fd_sc_hd__mux2_1
XFILLER_220_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13531_ _05936_ _06164_ _06219_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__a21o_1
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10743_ rbzero.tex_g0\[58\] rbzero.tex_g0\[57\] _03593_ vssd1 vssd1 vccd1 vccd1 _03594_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16250_ _08859_ _08860_ vssd1 vssd1 vccd1 vccd1 _08861_ sky130_fd_sc_hd__xor2_1
X_13462_ _06060_ _06063_ _06064_ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__a21o_1
XFILLER_55_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10674_ rbzero.tex_g1\[26\] rbzero.tex_g1\[27\] _03552_ vssd1 vssd1 vccd1 vccd1 _03558_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15201_ _07814_ _07685_ vssd1 vssd1 vccd1 vccd1 _07815_ sky130_fd_sc_hd__nor2_1
XFILLER_139_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12413_ _05104_ _05105_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__nand2_1
XFILLER_107_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16181_ _04938_ rbzero.wall_tracer.stepDistX\[5\] vssd1 vssd1 vccd1 vccd1 _08793_
+ sky130_fd_sc_hd__nand2_2
XFILLER_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13393_ _06073_ _06074_ _06080_ _06081_ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__a31o_1
XFILLER_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15132_ _07380_ _07743_ _07744_ _07745_ vssd1 vssd1 vccd1 vccd1 _07746_ sky130_fd_sc_hd__a22oi_2
XFILLER_177_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12344_ _05030_ _05033_ _05036_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__or3b_1
XFILLER_193_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15063_ _07674_ _07676_ vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19940_ _03117_ vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__clkinv_2
XFILLER_182_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12275_ rbzero.wall_tracer.trackDistX\[-12\] vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__inv_2
XFILLER_141_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14014_ _06697_ _06702_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__or2_1
X_11226_ _03944_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__buf_4
XFILLER_141_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19871_ _03110_ vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__clkinv_2
XFILLER_218_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18822_ _03729_ _02540_ _02541_ _02197_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__a31o_1
XTAP_6150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11157_ rbzero.texV\[8\] _03875_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__xnor2_1
XTAP_6161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18753_ _02473_ _02474_ _02475_ _02476_ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__a211o_1
XTAP_5460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15965_ _08573_ _08575_ _08578_ vssd1 vssd1 vccd1 vccd1 _08579_ sky130_fd_sc_hd__a21oi_1
XFILLER_114_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11088_ _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__clkinv_2
XTAP_5471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17704_ _10130_ _10131_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__nor2_1
XFILLER_209_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14916_ _07523_ _07524_ _07529_ vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__or3_1
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18684_ rbzero.debug_overlay.vplaneY\[-6\] _02396_ vssd1 vssd1 vccd1 vccd1 _02413_
+ sky130_fd_sc_hd__nand2_1
XFILLER_97_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15896_ _07880_ vssd1 vssd1 vccd1 vccd1 _08510_ sky130_fd_sc_hd__clkbuf_4
XFILLER_188_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17635_ _10058_ _10170_ vssd1 vssd1 vccd1 vccd1 _10171_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14847_ rbzero.wall_tracer.visualWallDist\[-7\] _03795_ _04936_ vssd1 vssd1 vccd1
+ vccd1 _07461_ sky130_fd_sc_hd__a21oi_1
XFILLER_149_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17566_ _10101_ _10102_ vssd1 vssd1 vccd1 vccd1 _10103_ sky130_fd_sc_hd__xnor2_1
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14778_ _05113_ _07390_ _07391_ _07351_ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__o211a_1
XFILLER_223_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19305_ rbzero.pov.spi_counter\[1\] rbzero.pov.spi_counter\[0\] _02837_ vssd1 vssd1
+ vccd1 vccd1 _02840_ sky130_fd_sc_hd__and3_1
X_16517_ _09124_ _09125_ vssd1 vssd1 vccd1 vccd1 _09126_ sky130_fd_sc_hd__xnor2_1
XFILLER_205_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13729_ _06405_ _06417_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__xnor2_2
XFILLER_182_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17497_ _10030_ _10031_ _10032_ vssd1 vssd1 vccd1 vccd1 _10034_ sky130_fd_sc_hd__o21a_1
XFILLER_149_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19236_ _02800_ vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__clkbuf_1
X_16448_ _07847_ _08923_ vssd1 vssd1 vccd1 vccd1 _09058_ sky130_fd_sc_hd__nor2_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19167_ _09247_ _02758_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__and2_1
X_16379_ _08983_ _08988_ vssd1 vssd1 vccd1 vccd1 _08989_ sky130_fd_sc_hd__xnor2_1
XFILLER_192_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18118_ _01894_ _01898_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__xor2_1
XFILLER_195_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19098_ net44 rbzero.spi_registers.sclk_buffer\[0\] _02708_ vssd1 vssd1 vccd1 vccd1
+ _02713_ sky130_fd_sc_hd__mux2_1
XFILLER_133_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18049_ _01820_ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__inv_2
XFILLER_144_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21060_ _00109_ _01076_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20011_ _03123_ vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__clkinv_2
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20913_ net78 _00929_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20844_ _00062_ _00860_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_230_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20775_ net88 _00791_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout56 net57 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_2
Xfanout67 net69 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_2
XFILLER_211_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout78 net1 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_202_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout89 net98 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10390_ rbzero.tex_r1\[31\] rbzero.tex_r1\[32\] _03400_ vssd1 vssd1 vccd1 vccd1 _03407_
+ sky130_fd_sc_hd__mux2_1
XFILLER_164_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21327_ _00350_ _01343_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12060_ net21 vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__buf_2
XFILLER_123_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21258_ _00307_ _01274_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11011_ _03732_ _03734_ _03738_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__o21ai_1
X_20209_ _03221_ _03224_ _03222_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__a21boi_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21189_ _00238_ _01205_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_237_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15750_ _08360_ _08363_ vssd1 vssd1 vccd1 vccd1 _08364_ sky130_fd_sc_hd__xor2_1
X_12962_ _05626_ _05630_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__nand2_2
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14701_ rbzero.wall_tracer.stepDistX\[5\] _07221_ _07316_ vssd1 vssd1 vccd1 vccd1
+ _07325_ sky130_fd_sc_hd__mux2_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ net10 net11 net12 vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__a21o_1
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _05576_ _05581_ _05538_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__mux2_1
X_15681_ _07481_ _07482_ vssd1 vssd1 vccd1 vccd1 _08295_ sky130_fd_sc_hd__and2_1
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17420_ _09956_ _09957_ vssd1 vssd1 vccd1 vccd1 _09958_ sky130_fd_sc_hd__nand2_1
XFILLER_2_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.trackDistY\[1\] _07258_
+ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__mux2_1
X_11844_ rbzero.tex_b1\[23\] rbzero.tex_b1\[22\] _04544_ vssd1 vssd1 vccd1 vccd1 _04558_
+ sky130_fd_sc_hd__mux2_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ rbzero.wall_tracer.trackDistX\[3\] rbzero.wall_tracer.stepDistX\[3\] vssd1
+ vssd1 vccd1 vccd1 _09890_ sky130_fd_sc_hd__or2_1
X_14563_ _05401_ _06988_ _05406_ _06985_ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__a211o_1
XFILLER_18_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ rbzero.tex_b0\[19\] rbzero.tex_b0\[18\] _04001_ vssd1 vssd1 vccd1 vccd1 _04490_
+ sky130_fd_sc_hd__mux2_1
XFILLER_246_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _08910_ _08911_ _08904_ vssd1 vssd1 vccd1 vccd1 _08913_ sky130_fd_sc_hd__a21oi_1
XFILLER_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13514_ _06201_ _06202_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__nor2_1
X_10726_ rbzero.tex_g1\[1\] rbzero.tex_g1\[2\] _03299_ vssd1 vssd1 vccd1 vccd1 _03585_
+ sky130_fd_sc_hd__mux2_1
X_17282_ _09818_ _09819_ vssd1 vssd1 vccd1 vccd1 _09821_ sky130_fd_sc_hd__and2_1
XFILLER_201_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14494_ _07176_ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__buf_2
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19021_ _02671_ vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__clkbuf_1
X_16233_ _08841_ _08843_ vssd1 vssd1 vccd1 vccd1 _08844_ sky130_fd_sc_hd__nor2_2
X_13445_ _06127_ _06128_ _06129_ _06131_ _06133_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__a32o_1
XFILLER_16_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10657_ rbzero.tex_g1\[34\] rbzero.tex_g1\[35\] _03541_ vssd1 vssd1 vccd1 vccd1 _03549_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16164_ _08774_ _08775_ vssd1 vssd1 vccd1 vccd1 _08776_ sky130_fd_sc_hd__xor2_1
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13376_ _06060_ _06063_ _06064_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__a21oi_1
XFILLER_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10588_ rbzero.tex_r0\[4\] rbzero.tex_r0\[3\] _03512_ vssd1 vssd1 vccd1 vccd1 _03513_
+ sky130_fd_sc_hd__mux2_1
X_12327_ rbzero.wall_tracer.trackDistX\[-9\] _05020_ rbzero.wall_tracer.trackDistY\[-12\]
+ _04969_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__a22o_1
X_15115_ _03794_ rbzero.wall_tracer.stepDistY\[-2\] vssd1 vssd1 vccd1 vccd1 _07729_
+ sky130_fd_sc_hd__nor2_1
XFILLER_138_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16095_ _08585_ _08706_ _04933_ vssd1 vssd1 vccd1 vccd1 _08708_ sky130_fd_sc_hd__a21o_1
XFILLER_127_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15046_ _07342_ _05073_ _07659_ _07337_ vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__o211a_1
XFILLER_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19923_ _03115_ vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__clkinv_2
X_12258_ _04949_ _04951_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__nand2_1
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11209_ _03914_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__clkbuf_4
XFILLER_110_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19854_ _03108_ vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__clkinv_2
XFILLER_190_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12189_ net38 vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__inv_2
XFILLER_214_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18805_ _02524_ _02525_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__xnor2_1
XFILLER_205_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19785_ _09247_ _03088_ _03089_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__and3_1
XFILLER_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16997_ _09536_ _09537_ vssd1 vssd1 vccd1 vccd1 _09538_ sky130_fd_sc_hd__nand2_1
XFILLER_83_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18736_ _04260_ rbzero.debug_overlay.vplaneY\[-6\] vssd1 vssd1 vccd1 vccd1 _02461_
+ sky130_fd_sc_hd__or2_1
X_15948_ _08460_ _08560_ vssd1 vssd1 vccd1 vccd1 _08562_ sky130_fd_sc_hd__or2_1
XTAP_5290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18667_ rbzero.debug_overlay.vplaneY\[-7\] _02393_ vssd1 vssd1 vccd1 vccd1 _02397_
+ sky130_fd_sc_hd__nand2_1
XFILLER_97_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15879_ _08483_ _08491_ _08492_ vssd1 vssd1 vccd1 vccd1 _08493_ sky130_fd_sc_hd__nand3_1
XFILLER_52_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17618_ _10051_ _10054_ _10052_ vssd1 vssd1 vccd1 vccd1 _10154_ sky130_fd_sc_hd__a21boi_1
X_18598_ _02275_ rbzero.wall_tracer.rayAddendX\[10\] vssd1 vssd1 vccd1 vccd1 _02337_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_149_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17549_ _10070_ _10085_ vssd1 vssd1 vccd1 vccd1 _10086_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20560_ net130 _00576_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19219_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.new_sky\[4\] _02786_
+ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__mux2_1
XFILLER_192_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20491_ net114 _00507_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_180_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21112_ _00161_ _01128_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21043_ _00092_ _01059_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20827_ _00045_ _00843_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_243_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11560_ _04229_ _04241_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__nor2_1
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20758_ net106 _00774_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_sky sky130_fd_sc_hd__dfxtp_1
XFILLER_211_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10511_ _03472_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11491_ _04201_ _04208_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__nor2_2
XFILLER_17_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20689_ net71 _00705_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[69\] sky130_fd_sc_hd__dfxtp_1
XFILLER_183_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13230_ _05887_ _05888_ _05615_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a21oi_1
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10442_ _03434_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13161_ _05624_ _05746_ _05749_ _05621_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__o22a_1
XFILLER_137_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10373_ rbzero.tex_r1\[39\] rbzero.tex_r1\[40\] _03389_ vssd1 vssd1 vccd1 vccd1 _03398_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12112_ _04778_ _04796_ _04818_ _04819_ vssd1 vssd1 vccd1 vccd1 o_gpout[3] sky130_fd_sc_hd__o31a_4
XFILLER_163_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13092_ _05737_ _05780_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16920_ _08787_ _09207_ vssd1 vssd1 vccd1 vccd1 _09462_ sky130_fd_sc_hd__and2_1
X_12043_ _04747_ _04751_ _04721_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__o21ba_1
XFILLER_219_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16851_ _08592_ _08717_ _08855_ _08507_ vssd1 vssd1 vccd1 vccd1 _09393_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_120_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15802_ _08413_ _08415_ vssd1 vssd1 vccd1 vccd1 _08416_ sky130_fd_sc_hd__nor2_1
XFILLER_65_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19570_ rbzero.pov.ready _02834_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__and2_2
X_16782_ _09303_ _09328_ _09329_ _09282_ vssd1 vssd1 vccd1 vccd1 _09330_ sky130_fd_sc_hd__a31o_1
XFILLER_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13994_ _06636_ _06638_ _06657_ _06682_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__a31o_1
XFILLER_150_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18521_ _02241_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__inv_2
XFILLER_98_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15733_ _08343_ _08345_ _08346_ vssd1 vssd1 vccd1 vccd1 _08347_ sky130_fd_sc_hd__a21o_1
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12945_ _05526_ _05546_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__nand2_4
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18452_ rbzero.wall_tracer.rayAddendX\[-1\] _02197_ _02201_ _02157_ vssd1 vssd1 vccd1
+ vccd1 _02202_ sky130_fd_sc_hd__a22o_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15664_ _08273_ _08276_ _08277_ vssd1 vssd1 vccd1 vccd1 _08278_ sky130_fd_sc_hd__o21a_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _05564_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__inv_2
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17403_ _09933_ _09940_ vssd1 vssd1 vccd1 vccd1 _09941_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14615_ _07245_ _07271_ _07272_ _07251_ vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__o211a_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _07332_ _02138_ _02039_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__o21a_1
XFILLER_159_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11827_ rbzero.tex_b1\[40\] _04119_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__and2_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15595_ _08194_ _08208_ vssd1 vssd1 vccd1 vccd1 _08209_ sky130_fd_sc_hd__xor2_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17334_ _09870_ _09872_ vssd1 vssd1 vccd1 vccd1 _09873_ sky130_fd_sc_hd__xor2_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14546_ _07218_ vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__clkbuf_1
X_11758_ rbzero.tex_b0\[37\] rbzero.tex_b0\[36\] _03904_ vssd1 vssd1 vccd1 vccd1 _04473_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10709_ _03576_ vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__clkbuf_1
X_17265_ _09802_ _09803_ vssd1 vssd1 vccd1 vccd1 _09804_ sky130_fd_sc_hd__nor2_1
XFILLER_144_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14477_ _07130_ _07108_ vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__nand2_2
XFILLER_174_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11689_ rbzero.tex_g1\[10\] _03959_ _03916_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__a21o_1
X_19004_ rbzero.pov.spi_buffer\[49\] rbzero.pov.ready_buffer\[49\] _02662_ vssd1 vssd1
+ vccd1 vccd1 _02663_ sky130_fd_sc_hd__mux2_1
XFILLER_128_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16216_ _08710_ _08827_ vssd1 vssd1 vccd1 vccd1 _08828_ sky130_fd_sc_hd__xnor2_4
X_13428_ _06102_ _06104_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__and2_1
XFILLER_31_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17196_ _09733_ _09735_ vssd1 vssd1 vccd1 vccd1 _09736_ sky130_fd_sc_hd__nand2_1
XFILLER_155_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16147_ _08757_ _08758_ vssd1 vssd1 vccd1 vccd1 _08759_ sky130_fd_sc_hd__xnor2_1
X_13359_ _06003_ _06004_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__xnor2_1
XFILLER_142_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16078_ _08689_ _08690_ vssd1 vssd1 vccd1 vccd1 _08691_ sky130_fd_sc_hd__nand2_1
XFILLER_29_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15029_ rbzero.debug_overlay.playerY\[-9\] _03793_ _04927_ _07642_ vssd1 vssd1 vccd1
+ vccd1 _07643_ sky130_fd_sc_hd__o211a_1
X_19906_ _03113_ vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__clkinv_2
XFILLER_123_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19837_ _02862_ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__buf_4
XFILLER_111_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19768_ _04110_ _04106_ _04114_ _03076_ _04920_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__o41a_1
Xinput2 i_debug_vec_overlay vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_4
XFILLER_216_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18719_ _02427_ _02430_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__or2_1
XFILLER_232_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19699_ rbzero.debug_overlay.playerY\[5\] _03050_ _03053_ _03012_ vssd1 vssd1 vccd1
+ vccd1 _03054_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20612_ net92 _00628_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20543_ net137 _00559_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20474_ net94 _00490_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_118_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21026_ net93 _01042_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10991_ rbzero.tex_b0\[4\] rbzero.tex_b0\[3\] _03715_ vssd1 vssd1 vccd1 vccd1 _03724_
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12730_ _05417_ _05418_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__nand2_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12661_ _05337_ _05349_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__xnor2_4
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14400_ _05569_ _07088_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__or2_1
X_11612_ rbzero.tex_g0\[13\] rbzero.tex_g0\[12\] _04148_ vssd1 vssd1 vccd1 vccd1 _04329_
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15380_ _07992_ _07993_ vssd1 vssd1 vccd1 vccd1 _07994_ sky130_fd_sc_hd__and2_1
X_12592_ _05220_ _05279_ _05280_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__a21o_1
XFILLER_180_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14331_ _07019_ _06969_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11543_ rbzero.debug_overlay.vplaneY\[-4\] _04242_ _04245_ _04260_ vssd1 vssd1 vccd1
+ vccd1 _04261_ sky130_fd_sc_hd__a22o_1
XFILLER_184_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17050_ _09463_ _09461_ _09467_ _09465_ vssd1 vssd1 vccd1 vccd1 _09591_ sky130_fd_sc_hd__o31ai_1
X_14262_ _06940_ _06942_ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__nand2_1
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11474_ _03896_ _04135_ _04157_ _04174_ _04191_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__o32a_1
X_16001_ _08590_ _08613_ vssd1 vssd1 vccd1 vccd1 _08614_ sky130_fd_sc_hd__xnor2_1
XFILLER_171_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13213_ _05885_ _05901_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__xor2_1
XFILLER_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10425_ _03425_ vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14193_ _06691_ _06881_ vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__xor2_1
XFILLER_124_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13144_ _05698_ _05735_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__xor2_1
XFILLER_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10356_ _03388_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__clkbuf_4
XFILLER_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17952_ _01640_ _01641_ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__nor2_1
XFILLER_174_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13075_ _05620_ _05649_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__and2b_1
XFILLER_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10287_ _03352_ vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_238_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16903_ _09443_ _09444_ vssd1 vssd1 vccd1 vccd1 _09445_ sky130_fd_sc_hd__nand2_1
X_12026_ net6 vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__inv_2
XFILLER_111_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17883_ _01656_ _01665_ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__nand2_1
XFILLER_238_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19622_ rbzero.debug_overlay.playerX\[3\] _02991_ vssd1 vssd1 vccd1 vccd1 _02994_
+ sky130_fd_sc_hd__and2_1
XFILLER_120_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16834_ _09135_ _09138_ _09375_ vssd1 vssd1 vccd1 vccd1 _09376_ sky130_fd_sc_hd__a21oi_2
XFILLER_66_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19553_ _02945_ vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16765_ _09311_ _09312_ _09313_ vssd1 vssd1 vccd1 vccd1 _09315_ sky130_fd_sc_hd__o21ai_1
XFILLER_150_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13977_ _06612_ _06611_ _06516_ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__a21o_1
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18504_ _02245_ _02246_ _02248_ _02249_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__o211ai_2
X_15716_ _08324_ _08328_ _08329_ _08289_ vssd1 vssd1 vccd1 vccd1 _08330_ sky130_fd_sc_hd__a211oi_2
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12928_ _05613_ _05614_ _05616_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__or3_1
X_19484_ _02909_ vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__clkbuf_1
X_16696_ rbzero.traced_texa\[-1\] _09264_ _09263_ rbzero.wall_tracer.visualWallDist\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__a22o_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18435_ _03730_ _02185_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__nor2_1
XFILLER_221_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15647_ _08252_ _08259_ vssd1 vssd1 vccd1 vccd1 _08261_ sky130_fd_sc_hd__nor2_1
XFILLER_59_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12859_ _05539_ _05547_ _05501_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__mux2_1
XFILLER_146_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18366_ _04992_ _02001_ _02124_ vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__a21oi_1
X_15578_ _08130_ _08145_ vssd1 vssd1 vccd1 vccd1 _08192_ sky130_fd_sc_hd__xnor2_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17317_ _09849_ _09855_ vssd1 vssd1 vccd1 vccd1 _09856_ sky130_fd_sc_hd__xor2_1
XFILLER_119_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14529_ _07177_ _07169_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__or2_1
X_18297_ _04953_ _07702_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__nor2_1
XFILLER_119_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17248_ _09785_ _09786_ vssd1 vssd1 vccd1 vccd1 _09787_ sky130_fd_sc_hd__nor2_1
XFILLER_174_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17179_ _07814_ _09463_ _09467_ _09603_ _09465_ vssd1 vssd1 vccd1 vccd1 _09719_ sky130_fd_sc_hd__o41a_1
XFILLER_116_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20190_ _03206_ _03210_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__nand2_1
XFILLER_118_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_40 rbzero.wall_tracer.visualWallDist\[-9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20526_ net123 _00542_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20457_ net94 _00007_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10210_ _03312_ vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11190_ _03908_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__buf_4
X_20388_ net135 _00419_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_175_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13900_ _06510_ _06586_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__nor2_1
XFILLER_48_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21009_ net80 _01025_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-7\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_5867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14880_ rbzero.debug_overlay.playerX\[-1\] vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__inv_2
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13831_ _06468_ _06473_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__xor2_1
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16550_ _09121_ _09158_ vssd1 vssd1 vccd1 vccd1 _09159_ sky130_fd_sc_hd__xnor2_1
XFILLER_1_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13762_ _06372_ _06399_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__nand2_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10974_ _03444_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__clkbuf_4
XFILLER_21_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15501_ _08097_ _08098_ vssd1 vssd1 vccd1 vccd1 _08115_ sky130_fd_sc_hd__xnor2_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12713_ _05310_ _05322_ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__and2_1
XFILLER_56_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16481_ _09089_ _09090_ vssd1 vssd1 vccd1 vccd1 _09091_ sky130_fd_sc_hd__nor2_1
XFILLER_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13693_ _06348_ _06381_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__and2_1
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18220_ rbzero.wall_tracer.trackDistY\[-12\] rbzero.wall_tracer.stepDistY\[-12\]
+ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__or2_1
X_15432_ _04936_ _07362_ _07363_ _07376_ vssd1 vssd1 vccd1 vccd1 _08046_ sky130_fd_sc_hd__o31a_4
XFILLER_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12644_ _05295_ _05265_ _05270_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__and3_1
X_18151_ _01927_ _01930_ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__xnor2_1
XFILLER_180_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15363_ _07976_ _07486_ vssd1 vssd1 vccd1 vccd1 _07977_ sky130_fd_sc_hd__xnor2_1
X_12575_ _05227_ _05229_ _05233_ _05263_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__a211o_1
XFILLER_129_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17102_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.stepDistX\[1\] vssd1
+ vssd1 vccd1 vccd1 _09643_ sky130_fd_sc_hd__nand2_1
XFILLER_156_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14314_ _06997_ _07002_ vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__or2_1
XFILLER_184_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18082_ _01768_ _01862_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__xnor2_1
X_11526_ _04225_ _04208_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__nor2_4
XFILLER_117_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15294_ _07810_ _07787_ vssd1 vssd1 vccd1 vccd1 _07908_ sky130_fd_sc_hd__or2b_1
XFILLER_102_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17033_ _07631_ _09429_ vssd1 vssd1 vccd1 vccd1 _09574_ sky130_fd_sc_hd__nor2_1
XFILLER_172_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14245_ _05959_ _06542_ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__or2_1
X_11457_ rbzero.tex_r1\[15\] rbzero.tex_r1\[14\] _04168_ vssd1 vssd1 vccd1 vccd1 _04175_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10408_ _03416_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__clkbuf_1
X_14176_ _06848_ _06864_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__nand2_1
XFILLER_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11388_ gpout0.hpos\[2\] _04085_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__nand2_1
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13127_ _05687_ _05695_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10339_ rbzero.tex_r1\[55\] rbzero.tex_r1\[56\] _03377_ vssd1 vssd1 vccd1 vccd1 _03380_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18984_ _02652_ vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__clkbuf_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17935_ _01716_ _01717_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__and2_1
X_13058_ _05621_ _05746_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__nor2_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12009_ net4 vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__buf_2
XFILLER_94_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17866_ _01547_ _01560_ _01559_ vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__a21o_1
XFILLER_152_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16817_ rbzero.wall_tracer.trackDistX\[-2\] _09301_ _09354_ _09360_ vssd1 vssd1 vccd1
+ vccd1 _00551_ sky130_fd_sc_hd__o22a_1
X_19605_ _02956_ _02979_ _02980_ _02978_ vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__o211a_1
XFILLER_113_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17797_ _01573_ _01580_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__xor2_1
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19536_ rbzero.pov.spi_buffer\[63\] rbzero.pov.spi_buffer\[64\] _02932_ vssd1 vssd1
+ vccd1 vccd1 _02937_ sky130_fd_sc_hd__mux2_1
XFILLER_59_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16748_ _09279_ _09298_ _09299_ _09283_ vssd1 vssd1 vccd1 vccd1 _09300_ sky130_fd_sc_hd__a31o_1
XFILLER_81_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19467_ rbzero.pov.spi_buffer\[30\] rbzero.pov.spi_buffer\[31\] _02899_ vssd1 vssd1
+ vccd1 vccd1 _02901_ sky130_fd_sc_hd__mux2_1
X_16679_ rbzero.row_render.texu\[3\] _09260_ _09258_ rbzero.wall_tracer.texu\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__a22o_1
XFILLER_185_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18418_ rbzero.debug_overlay.vplaneX\[-7\] _02168_ vssd1 vssd1 vccd1 vccd1 _02170_
+ sky130_fd_sc_hd__or2_1
XFILLER_179_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19398_ _02863_ vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__clkinv_2
XFILLER_210_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18349_ _02107_ _02108_ _02109_ vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__or3_1
XFILLER_163_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21360_ _00383_ _01376_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20311_ rbzero.traced_texVinit\[2\] _09266_ _08564_ _09261_ vssd1 vssd1 vccd1 vccd1
+ _01396_ sky130_fd_sc_hd__a22o_1
XFILLER_198_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21291_ net134 _01307_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20242_ _03253_ vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__clkinv_2
XFILLER_200_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20173_ _03093_ _03196_ _03198_ _03064_ rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1
+ _01318_ sky130_fd_sc_hd__a32o_1
XFILLER_143_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10690_ _03566_ vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12360_ rbzero.debug_overlay.facingY\[-1\] rbzero.wall_tracer.rayAddendY\[7\] vssd1
+ vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__nand2_1
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11311_ gpout0.hpos\[9\] _04029_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__nor2_4
X_20509_ net129 _00525_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-2\] sky130_fd_sc_hd__dfxtp_1
X_12291_ rbzero.wall_tracer.trackDistX\[3\] vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__inv_2
XFILLER_154_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14030_ _06101_ _06342_ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__nor2_1
XFILLER_180_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11242_ _03903_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__buf_4
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11173_ _03888_ _03890_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__or2_1
XTAP_7055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15981_ _08067_ vssd1 vssd1 vccd1 vccd1 _08594_ sky130_fd_sc_hd__clkbuf_4
XTAP_5620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17720_ _09345_ _01504_ vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__nand2_1
XTAP_6387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14932_ rbzero.debug_overlay.playerX\[-2\] _07492_ vssd1 vssd1 vccd1 vccd1 _07546_
+ sky130_fd_sc_hd__xnor2_1
XTAP_5664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17651_ _01434_ _01435_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__xnor2_1
XTAP_5697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ _07378_ _07387_ _07399_ _07424_ vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__o22ai_1
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16602_ _09209_ _09210_ vssd1 vssd1 vccd1 vccd1 _09211_ sky130_fd_sc_hd__xnor2_1
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13814_ _06457_ _06498_ _06502_ vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__o21a_1
XFILLER_169_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17582_ _10116_ _10117_ _10110_ vssd1 vssd1 vccd1 vccd1 _10119_ sky130_fd_sc_hd__a21o_1
XFILLER_235_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14794_ _07349_ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__clkbuf_4
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19321_ rbzero.pov.spi_counter\[5\] _02849_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__and2_1
X_16533_ _09017_ _09021_ vssd1 vssd1 vccd1 vccd1 _09142_ sky130_fd_sc_hd__nand2_1
XFILLER_216_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13745_ _06418_ _06433_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10957_ _03706_ vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19252_ _02809_ vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16464_ _08914_ _08940_ _09073_ vssd1 vssd1 vccd1 vccd1 _09074_ sky130_fd_sc_hd__a21bo_1
XFILLER_143_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13676_ _05722_ _06306_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__nor2_1
XFILLER_32_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10888_ rbzero.tex_b0\[53\] rbzero.tex_b0\[52\] _03660_ vssd1 vssd1 vccd1 vccd1 _03670_
+ sky130_fd_sc_hd__mux2_1
X_18203_ _01892_ _01900_ _01982_ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__a21oi_1
XFILLER_188_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15415_ _08002_ _08028_ vssd1 vssd1 vccd1 vccd1 _08029_ sky130_fd_sc_hd__nor2_1
XPHY_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12627_ _05199_ _05204_ _05271_ _05276_ _05296_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__o41a_2
X_19183_ rbzero.spi_registers.new_floor\[3\] rbzero.spi_registers.got_new_floor _02724_
+ _02753_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__a31o_1
XPHY_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16395_ _08863_ _08870_ _09004_ vssd1 vssd1 vccd1 vccd1 _09005_ sky130_fd_sc_hd__a21oi_1
XPHY_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18134_ _01913_ _01834_ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__and2b_1
XFILLER_200_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15346_ _07930_ _07959_ vssd1 vssd1 vccd1 vccd1 _07960_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12558_ _05149_ _05246_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__xnor2_2
XFILLER_129_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18065_ _01843_ _01845_ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__xnor2_1
X_11509_ _03783_ _04223_ _04213_ _04226_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__a211o_1
X_15277_ _07469_ _07890_ _07800_ _07388_ vssd1 vssd1 vccd1 vccd1 _07891_ sky130_fd_sc_hd__o22ai_1
XFILLER_184_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12489_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[9\] vssd1
+ vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__or2_1
XFILLER_67_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17016_ _09406_ _09411_ vssd1 vssd1 vccd1 vccd1 _09557_ sky130_fd_sc_hd__and2b_1
X_14228_ _06889_ _06914_ _06916_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__o21ba_1
XFILLER_160_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14159_ _06435_ _06542_ _06847_ vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__or3_1
XFILLER_125_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18967_ _02643_ vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__clkbuf_1
XFILLER_234_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17918_ _01518_ _01700_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__xnor2_1
XFILLER_239_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18898_ rbzero.pov.spi_done _03292_ vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__nand2_2
XFILLER_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17849_ _01630_ _01631_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__nand2_1
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20860_ _00078_ _00876_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19519_ rbzero.pov.spi_buffer\[55\] rbzero.pov.spi_buffer\[56\] _02921_ vssd1 vssd1
+ vccd1 vccd1 _02928_ sky130_fd_sc_hd__mux2_1
X_20791_ net91 _00807_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready sky130_fd_sc_hd__dfxtp_1
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21343_ _00366_ _01359_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21274_ _00323_ _01290_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20225_ _03234_ _03238_ _03235_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__o21ai_1
XFILLER_104_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20156_ _03182_ _03183_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__or2_1
XFILLER_58_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20087_ _03131_ vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__clkinv_2
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11860_ rbzero.tex_b1\[11\] _03938_ _03940_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__and3_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10811_ rbzero.tex_g0\[26\] rbzero.tex_g0\[25\] _03627_ vssd1 vssd1 vccd1 vccd1 _03630_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11791_ rbzero.tex_b0\[15\] rbzero.tex_b0\[14\] _03925_ vssd1 vssd1 vccd1 vccd1 _04506_
+ sky130_fd_sc_hd__mux2_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20989_ net65 _01005_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13530_ _05879_ _05935_ vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__and2_1
XFILLER_242_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10742_ _03445_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__clkbuf_4
XFILLER_246_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13461_ _06026_ _06065_ _06149_ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__or3b_1
X_10673_ _03557_ vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15200_ _07468_ vssd1 vssd1 vccd1 vccd1 _07814_ sky130_fd_sc_hd__clkbuf_4
X_12412_ _05061_ _05103_ _05059_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__a21o_1
X_16180_ _08790_ _08791_ vssd1 vssd1 vccd1 vccd1 _08792_ sky130_fd_sc_hd__and2_1
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13392_ _06075_ _06079_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__and2b_1
XFILLER_142_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15131_ _07388_ _07416_ vssd1 vssd1 vccd1 vccd1 _07745_ sky130_fd_sc_hd__nor2_1
XFILLER_139_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12343_ _05034_ _05035_ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__nor2_1
XFILLER_177_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15062_ _07455_ _07675_ vssd1 vssd1 vccd1 vccd1 _07676_ sky130_fd_sc_hd__nor2_1
X_12274_ rbzero.wall_tracer.trackDistX\[-11\] vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__inv_2
XFILLER_138_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14013_ _06651_ _06698_ _06699_ _06701_ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__o2bb2a_1
X_11225_ _03864_ _03894_ _03918_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__or3_4
XFILLER_175_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19870_ _02862_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__buf_4
X_11156_ _03873_ _03874_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__nor2_1
X_18821_ _02523_ _02534_ _02539_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__a21o_1
XTAP_6140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18752_ _02446_ _02457_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__nor2_1
XTAP_5450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15964_ _08576_ _08577_ vssd1 vssd1 vccd1 vccd1 _08578_ sky130_fd_sc_hd__nand2_1
X_11087_ _03801_ _03809_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__and2_1
XTAP_6195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17703_ _01448_ _01487_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__xnor2_1
XTAP_5472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14915_ _07349_ _07525_ _07526_ _07528_ _07352_ vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__a221o_4
XTAP_5494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18683_ _02157_ _02411_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__nor2_1
X_15895_ _08506_ _08508_ vssd1 vssd1 vccd1 vccd1 _08509_ sky130_fd_sc_hd__nand2_1
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17634_ _09571_ _08717_ vssd1 vssd1 vccd1 vccd1 _10170_ sky130_fd_sc_hd__nor2_1
XFILLER_188_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14846_ _07453_ _07459_ vssd1 vssd1 vccd1 vccd1 _07460_ sky130_fd_sc_hd__nand2_1
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17565_ _08760_ _09451_ vssd1 vssd1 vccd1 vccd1 _10102_ sky130_fd_sc_hd__nor2_1
XFILLER_205_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14777_ _07389_ _05113_ vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__nand2_1
XFILLER_51_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11989_ net52 _04664_ _04665_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__and3_1
XFILLER_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19304_ rbzero.pov.spi_counter\[0\] _02837_ _02839_ vssd1 vssd1 vccd1 vccd1 _00808_
+ sky130_fd_sc_hd__a21oi_1
X_16516_ _07515_ _08850_ vssd1 vssd1 vccd1 vccd1 _09125_ sky130_fd_sc_hd__nor2_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13728_ _06410_ _06415_ _06416_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__o21a_1
XFILLER_225_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17496_ _10030_ _10031_ _10032_ vssd1 vssd1 vccd1 vccd1 _10033_ sky130_fd_sc_hd__nor3_1
XFILLER_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19235_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.new_floor\[4\]
+ _02795_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__mux2_1
X_16447_ _07680_ _08787_ _09055_ _07838_ vssd1 vssd1 vccd1 vccd1 _09057_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_177_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13659_ _06339_ _06347_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__or2_1
XFILLER_20_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19166_ rbzero.spi_registers.new_sky\[3\] rbzero.color_sky\[3\] _02752_ vssd1 vssd1
+ vccd1 vccd1 _02758_ sky130_fd_sc_hd__mux2_1
X_16378_ _08986_ _08987_ vssd1 vssd1 vccd1 vccd1 _08988_ sky130_fd_sc_hd__and2b_1
XFILLER_192_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18117_ _01896_ _01897_ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__and2_1
XFILLER_30_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15329_ _07762_ _07934_ _07941_ vssd1 vssd1 vccd1 vccd1 _07943_ sky130_fd_sc_hd__a21o_1
XFILLER_121_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19097_ _02712_ vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18048_ _01823_ _01829_ rbzero.wall_tracer.trackDistX\[9\] _09276_ vssd1 vssd1 vccd1
+ vccd1 _00562_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_201_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20010_ _03123_ vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__clkinv_2
XFILLER_236_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19999_ _03122_ vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__clkinv_2
XFILLER_101_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20912_ net78 _00928_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_215_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ _00061_ _00859_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20774_ net102 _00790_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_223_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout57 net58 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_2
XFILLER_195_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout68 net69 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout79 net80 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__buf_2
XFILLER_91_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21326_ _00349_ _01342_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21257_ _00306_ _01273_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _03735_ _03737_ _03733_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__or3b_1
X_20208_ _03226_ _03227_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__and2b_1
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21188_ _00237_ _01204_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20139_ _03168_ _03169_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__xnor2_1
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ _05620_ _05649_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _07324_ vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__clkbuf_1
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ net12 net11 vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__nor2_1
XFILLER_85_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15680_ _07507_ _07645_ _08293_ _07882_ vssd1 vssd1 vccd1 vccd1 _08294_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12892_ _05577_ _05500_ _05579_ _05580_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__o211a_1
XFILLER_2_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14631_ _07245_ _07282_ _07283_ _07251_ vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__o211a_1
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11843_ rbzero.tex_b1\[21\] rbzero.tex_b1\[20\] _04544_ vssd1 vssd1 vccd1 vccd1 _04557_
+ sky130_fd_sc_hd__mux2_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17350_ rbzero.wall_tracer.trackDistX\[3\] rbzero.wall_tracer.stepDistX\[3\] vssd1
+ vssd1 vccd1 vccd1 _09889_ sky130_fd_sc_hd__nand2_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14562_ _07057_ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__inv_2
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _03994_ _04484_ _04488_ _03956_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__a211o_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _08904_ _08910_ _08911_ vssd1 vssd1 vccd1 vccd1 _08912_ sky130_fd_sc_hd__and3_1
XFILLER_201_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13513_ _05553_ _05701_ _06200_ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__a21oi_1
X_17281_ _09818_ _09819_ vssd1 vssd1 vccd1 vccd1 _09820_ sky130_fd_sc_hd__nor2_1
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ _03584_ vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__clkbuf_1
X_14493_ _05602_ _05577_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__or2_1
X_19020_ rbzero.pov.spi_buffer\[57\] rbzero.pov.ready_buffer\[57\] _02662_ vssd1 vssd1
+ vccd1 vccd1 _02671_ sky130_fd_sc_hd__mux2_1
X_16232_ _08715_ _08744_ _08842_ vssd1 vssd1 vccd1 vccd1 _08843_ sky130_fd_sc_hd__a21boi_1
XFILLER_186_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13444_ _06123_ _06132_ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__and2_1
XFILLER_146_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10656_ _03548_ vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16163_ _07858_ _07685_ vssd1 vssd1 vccd1 vccd1 _08775_ sky130_fd_sc_hd__nor2_1
X_13375_ _05992_ _06020_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__xnor2_1
X_10587_ _03445_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__clkbuf_4
XFILLER_154_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15114_ _07725_ _07727_ vssd1 vssd1 vccd1 vccd1 _07728_ sky130_fd_sc_hd__nand2_1
XFILLER_177_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12326_ rbzero.wall_tracer.trackDistY\[-9\] vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__inv_2
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16094_ _08585_ _08706_ vssd1 vssd1 vccd1 vccd1 _08707_ sky130_fd_sc_hd__nor2_1
XFILLER_182_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15045_ _07342_ _05196_ vssd1 vssd1 vccd1 vccd1 _07659_ sky130_fd_sc_hd__nand2_1
XFILLER_141_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19922_ _03115_ vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__clkinv_2
X_12257_ _04950_ rbzero.wall_tracer.trackDistY\[-2\] _04947_ rbzero.wall_tracer.trackDistY\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__o22a_1
XFILLER_218_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11208_ rbzero.tex_r0\[61\] rbzero.tex_r0\[60\] _03925_ vssd1 vssd1 vccd1 vccd1 _03927_
+ sky130_fd_sc_hd__mux2_1
X_12188_ _04883_ o_rgb[7] _04893_ net37 vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a211o_1
X_19853_ _03108_ vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__clkinv_2
XFILLER_229_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18804_ _02500_ _02503_ _02501_ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__o21bai_1
X_11139_ rbzero.traced_texVinit\[2\] rbzero.texV\[2\] _03857_ vssd1 vssd1 vccd1 vccd1
+ _03858_ sky130_fd_sc_hd__o21ai_2
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16996_ _08274_ _08596_ _08718_ _08985_ vssd1 vssd1 vccd1 vccd1 _09537_ sky130_fd_sc_hd__or4_1
X_19784_ _04632_ _04631_ _04628_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__a21o_1
XFILLER_205_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15947_ _08460_ _08560_ vssd1 vssd1 vccd1 vccd1 _08561_ sky130_fd_sc_hd__nand2_1
XFILLER_114_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18735_ _04260_ rbzero.debug_overlay.vplaneY\[-6\] vssd1 vssd1 vccd1 vccd1 _02460_
+ sky130_fd_sc_hd__nand2_1
XTAP_5280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18666_ rbzero.debug_overlay.vplaneY\[-7\] _02393_ vssd1 vssd1 vccd1 vccd1 _02396_
+ sky130_fd_sc_hd__or2_1
X_15878_ _08488_ _08489_ _08490_ vssd1 vssd1 vccd1 vccd1 _08492_ sky130_fd_sc_hd__a21o_1
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17617_ _10089_ _10048_ vssd1 vssd1 vccd1 vccd1 _10153_ sky130_fd_sc_hd__or2b_1
XFILLER_221_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14829_ rbzero.wall_tracer.visualWallDist\[-12\] _03795_ vssd1 vssd1 vccd1 vccd1
+ _07443_ sky130_fd_sc_hd__nand2_2
XFILLER_92_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18597_ _02191_ _02312_ _03729_ _02335_ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__o211a_1
XFILLER_240_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17548_ _10083_ _10084_ vssd1 vssd1 vccd1 vccd1 _10085_ sky130_fd_sc_hd__nor2_1
XFILLER_196_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17479_ _09878_ _09880_ _10016_ vssd1 vssd1 vccd1 vccd1 _10017_ sky130_fd_sc_hd__o21a_1
XFILLER_220_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19218_ _02790_ vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__clkbuf_1
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20490_ net112 _00506_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19149_ rbzero.spi_registers.new_leak\[2\] _02745_ vssd1 vssd1 vccd1 vccd1 _02748_
+ sky130_fd_sc_hd__or2_1
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21111_ _00160_ _01127_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21042_ _00091_ _01058_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_232_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20826_ _00044_ _00842_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20757_ net105 _00773_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10510_ rbzero.tex_r0\[41\] rbzero.tex_r0\[40\] _03468_ vssd1 vssd1 vccd1 vccd1 _03472_
+ sky130_fd_sc_hd__mux2_1
XFILLER_195_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11490_ _04203_ _04207_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__nand2_2
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20688_ net70 _00704_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[68\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10441_ rbzero.tex_r1\[7\] rbzero.tex_r1\[8\] _03433_ vssd1 vssd1 vccd1 vccd1 _03434_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13160_ _05747_ _05848_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__and2_1
XFILLER_152_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10372_ _03397_ vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12111_ o_rgb[7] _04779_ _04803_ _04809_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__nand4b_1
X_13091_ _05761_ _05779_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__xnor2_1
X_21309_ net114 _01325_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12042_ _04702_ _04748_ _04749_ gpout0.clk_div\[0\] _04750_ vssd1 vssd1 vccd1 vccd1
+ _04751_ sky130_fd_sc_hd__a221o_1
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16850_ _08592_ _08296_ _08716_ _08984_ vssd1 vssd1 vccd1 vccd1 _09392_ sky130_fd_sc_hd__or4_1
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15801_ _08356_ _08414_ vssd1 vssd1 vccd1 vccd1 _08415_ sky130_fd_sc_hd__nand2_1
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16781_ _09325_ _09326_ _09327_ vssd1 vssd1 vccd1 vccd1 _09329_ sky130_fd_sc_hd__o21ai_1
XFILLER_111_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13993_ _06641_ _06656_ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__nor2_1
XFILLER_115_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18520_ _02263_ _02264_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__nand2_1
XFILLER_219_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15732_ _08332_ _08342_ vssd1 vssd1 vccd1 vccd1 _08346_ sky130_fd_sc_hd__and2b_1
XFILLER_65_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ _05623_ _05632_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _02188_ _02200_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__xnor2_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ _08274_ _07971_ _08275_ vssd1 vssd1 vccd1 vccd1 _08277_ sky130_fd_sc_hd__or3_1
XFILLER_59_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12875_ _05556_ _05499_ _05558_ _05563_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__o211a_2
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17402_ _09934_ _09939_ vssd1 vssd1 vccd1 vccd1 _09940_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14614_ rbzero.wall_tracer.visualWallDist\[-5\] _07252_ vssd1 vssd1 vccd1 vccd1 _07272_
+ sky130_fd_sc_hd__or2_1
XFILLER_57_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _02136_ _02137_ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__xnor2_1
X_11826_ rbzero.tex_b1\[43\] rbzero.tex_b1\[42\] _03903_ vssd1 vssd1 vccd1 vccd1 _04540_
+ sky130_fd_sc_hd__mux2_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15594_ _08196_ _08206_ _08207_ vssd1 vssd1 vccd1 vccd1 _08208_ sky130_fd_sc_hd__a21oi_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17333_ _09717_ _09743_ _09871_ vssd1 vssd1 vccd1 vccd1 _09872_ sky130_fd_sc_hd__a21boi_1
XFILLER_226_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ rbzero.wall_tracer.stepDistY\[4\] _07217_ _07193_ vssd1 vssd1 vccd1 vccd1
+ _07218_ sky130_fd_sc_hd__mux2_1
XFILLER_159_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11757_ rbzero.tex_b0\[39\] rbzero.tex_b0\[38\] _03904_ vssd1 vssd1 vccd1 vccd1 _04472_
+ sky130_fd_sc_hd__mux2_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17264_ _08596_ _08725_ _09670_ _09669_ vssd1 vssd1 vccd1 vccd1 _09803_ sky130_fd_sc_hd__o31a_1
XFILLER_140_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10708_ rbzero.tex_g1\[10\] rbzero.tex_g1\[11\] _03574_ vssd1 vssd1 vccd1 vccd1 _03576_
+ sky130_fd_sc_hd__mux2_1
X_14476_ _07107_ _07106_ _07160_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__a21oi_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11688_ rbzero.tex_g1\[11\] _04143_ _04145_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__and3_1
XFILLER_179_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19003_ _02606_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__clkbuf_4
XFILLER_31_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16215_ _08825_ _08826_ vssd1 vssd1 vccd1 vccd1 _08827_ sky130_fd_sc_hd__and2_2
XFILLER_122_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13427_ _06028_ _06115_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__nand2_1
X_17195_ _09609_ _09732_ _09734_ _09476_ vssd1 vssd1 vccd1 vccd1 _09735_ sky130_fd_sc_hd__a211o_2
X_10639_ _03539_ vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16146_ _07742_ _07805_ vssd1 vssd1 vccd1 vccd1 _08758_ sky130_fd_sc_hd__or2_1
XFILLER_155_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13358_ _06002_ _06042_ _06043_ _06046_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__o22ai_2
XFILLER_128_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12309_ rbzero.wall_tracer.trackDistX\[5\] _05002_ _05001_ rbzero.wall_tracer.trackDistX\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__o22a_1
X_16077_ _08686_ _08688_ vssd1 vssd1 vccd1 vccd1 _08690_ sky130_fd_sc_hd__nand2_1
XFILLER_170_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13289_ _05937_ _05977_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__nor2_1
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15028_ rbzero.wall_tracer.visualWallDist\[-9\] rbzero.wall_tracer.state\[13\] vssd1
+ vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__or2_1
X_19905_ _03113_ vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__clkinv_2
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19836_ _03106_ vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__clkinv_2
XFILLER_233_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19767_ _04246_ _04632_ gpout0.vpos\[0\] _04628_ vssd1 vssd1 vccd1 vccd1 _03076_
+ sky130_fd_sc_hd__or4b_1
XFILLER_42_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput3 i_gpout0_sel[0] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_6
X_16979_ _09398_ _09401_ _09519_ vssd1 vssd1 vccd1 vccd1 _09520_ sky130_fd_sc_hd__a21oi_2
XFILLER_110_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18718_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__or2_1
X_19698_ rbzero.pov.ready_buffer\[58\] _02962_ _03052_ vssd1 vssd1 vccd1 vccd1 _03053_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_37_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18649_ rbzero.debug_overlay.vplaneY\[-6\] rbzero.wall_tracer.rayAddendY\[-6\] _02380_
+ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a21o_1
XFILLER_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20611_ net92 _00627_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_240_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20542_ net137 _00558_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20473_ net112 _00489_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_192_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21025_ net95 _01041_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10990_ _03723_ vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12660_ _05305_ _05336_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__nand2_1
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11611_ rbzero.tex_g0\[15\] rbzero.tex_g0\[14\] _04148_ vssd1 vssd1 vccd1 vccd1 _04328_
+ sky130_fd_sc_hd__mux2_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20809_ _00027_ _00825_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[10\] sky130_fd_sc_hd__dfxtp_1
X_12591_ _05143_ _05184_ _05185_ _05220_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__a211oi_4
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14330_ _06794_ _06966_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__nand2_1
XFILLER_204_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11542_ rbzero.debug_overlay.vplaneY\[-2\] vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__buf_2
XFILLER_195_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14261_ _06938_ _06940_ _06945_ _06949_ vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__and4_1
XFILLER_156_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11473_ _03985_ _04182_ _04190_ _04026_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__a31o_1
XFILLER_109_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16000_ _08591_ _08612_ vssd1 vssd1 vccd1 vccd1 _08613_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13212_ _05892_ _05899_ _05900_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__o21a_1
XFILLER_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10424_ rbzero.tex_r1\[15\] rbzero.tex_r1\[16\] _03422_ vssd1 vssd1 vccd1 vccd1 _03425_
+ sky130_fd_sc_hd__mux2_1
X_14192_ _05740_ _06542_ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__or2_1
XFILLER_178_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13143_ _05817_ _05830_ _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__a21o_1
XFILLER_152_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10355_ _03298_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__clkbuf_4
XFILLER_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17951_ _01732_ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__inv_2
X_13074_ _05648_ _05644_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__and2b_1
XFILLER_139_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ rbzero.tex_b1\[16\] rbzero.tex_b1\[17\] _03344_ vssd1 vssd1 vccd1 vccd1 _03352_
+ sky130_fd_sc_hd__mux2_1
XFILLER_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16902_ _09426_ _09194_ _09442_ vssd1 vssd1 vccd1 vccd1 _09444_ sky130_fd_sc_hd__nand3_1
X_12025_ net6 _04733_ _04718_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__o21ba_1
X_17882_ _01663_ _01664_ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__and2_1
XFILLER_238_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19621_ rbzero.debug_overlay.playerX\[2\] _02960_ _02993_ _02989_ vssd1 vssd1 vccd1
+ vccd1 _00971_ sky130_fd_sc_hd__a211o_1
X_16833_ _08429_ _09373_ _09126_ _09374_ vssd1 vssd1 vccd1 vccd1 _09375_ sky130_fd_sc_hd__o31a_1
XFILLER_226_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16764_ _09311_ _09312_ _09313_ vssd1 vssd1 vccd1 vccd1 _09314_ sky130_fd_sc_hd__or3_1
X_19552_ rbzero.pov.spi_buffer\[71\] rbzero.pov.spi_buffer\[72\] _02865_ vssd1 vssd1
+ vccd1 vccd1 _02945_ sky130_fd_sc_hd__mux2_1
X_13976_ _06516_ _06612_ _06611_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__nand3_1
XFILLER_47_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15715_ _08272_ _07986_ _08060_ _07400_ vssd1 vssd1 vccd1 vccd1 _08329_ sky130_fd_sc_hd__o22a_1
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18503_ _02247_ rbzero.wall_tracer.rayAddendX\[3\] vssd1 vssd1 vccd1 vccd1 _02249_
+ sky130_fd_sc_hd__or2_1
X_12927_ _05552_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__clkbuf_4
XFILLER_111_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16695_ rbzero.traced_texa\[-2\] _09264_ _09263_ rbzero.wall_tracer.visualWallDist\[-2\]
+ vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__a22o_1
X_19483_ rbzero.pov.spi_buffer\[38\] rbzero.pov.spi_buffer\[39\] _02899_ vssd1 vssd1
+ vccd1 vccd1 _02909_ sky130_fd_sc_hd__mux2_1
XFILLER_234_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15646_ _08252_ _08259_ vssd1 vssd1 vccd1 vccd1 _08260_ sky130_fd_sc_hd__xor2_1
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18434_ _02183_ _02184_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__xor2_1
X_12858_ _05372_ _05417_ _05463_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__mux2_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18365_ _09345_ _02123_ _01995_ _01721_ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__o211a_1
XFILLER_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11809_ rbzero.tex_b1\[55\] rbzero.tex_b1\[54\] _04032_ vssd1 vssd1 vccd1 vccd1 _04523_
+ sky130_fd_sc_hd__mux2_1
X_15577_ _08188_ _08190_ vssd1 vssd1 vccd1 vccd1 _08191_ sky130_fd_sc_hd__nor2_1
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12789_ _05477_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__buf_2
XFILLER_203_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _09850_ _09854_ vssd1 vssd1 vccd1 vccd1 _09855_ sky130_fd_sc_hd__xor2_1
XFILLER_175_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14528_ _07133_ _07074_ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__or2_1
XFILLER_187_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18296_ rbzero.wall_tracer.trackDistY\[-1\] rbzero.wall_tracer.stepDistY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__nor2_1
XFILLER_202_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17247_ _09777_ _09778_ _09784_ vssd1 vssd1 vccd1 vccd1 _09786_ sky130_fd_sc_hd__and3_1
XFILLER_179_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14459_ _05577_ _07140_ _07145_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__a21o_1
XFILLER_128_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17178_ _09592_ _09596_ vssd1 vssd1 vccd1 vccd1 _09718_ sky130_fd_sc_hd__nand2_1
XFILLER_157_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16129_ _08739_ _08740_ vssd1 vssd1 vccd1 vccd1 _08741_ sky130_fd_sc_hd__nor2_1
XFILLER_157_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19819_ _03105_ vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__clkinv_2
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_30 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_41 rbzero.wall_tracer.visualWallDist\[-9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20525_ net124 _00541_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20456_ net119 _00006_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20387_ net135 _00418_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_106_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21008_ net80 _01024_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_87_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13830_ _06512_ _06514_ _06518_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__a21boi_1
XFILLER_25_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13761_ _06404_ _06449_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__nor2_1
X_10973_ _03714_ vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15500_ _08113_ _08103_ vssd1 vssd1 vccd1 vccd1 _08114_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12712_ _05400_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__buf_4
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16480_ _09087_ _09088_ _08974_ vssd1 vssd1 vccd1 vccd1 _09090_ sky130_fd_sc_hd__a21oi_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13692_ _06339_ _06347_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__nand2_1
XFILLER_243_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15431_ _07964_ _07554_ vssd1 vssd1 vccd1 vccd1 _08045_ sky130_fd_sc_hd__nand2_1
X_12643_ _05296_ _05271_ _05330_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18150_ _01928_ _01929_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15362_ _07487_ _07477_ vssd1 vssd1 vccd1 vccd1 _07976_ sky130_fd_sc_hd__nand2_1
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12574_ _05237_ _05239_ _05262_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__a21o_1
XFILLER_184_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17101_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.stepDistX\[1\] vssd1
+ vssd1 vccd1 vccd1 _09642_ sky130_fd_sc_hd__or2_1
XFILLER_129_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14313_ _05593_ _07001_ vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__and2_1
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18081_ _10095_ _08718_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__nor2_1
XFILLER_141_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11525_ _04216_ _04208_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__nor2_2
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15293_ _07904_ _07905_ _07782_ _07813_ vssd1 vssd1 vccd1 vccd1 _07907_ sky130_fd_sc_hd__a211o_1
XFILLER_32_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17032_ _09570_ _09572_ vssd1 vssd1 vccd1 vccd1 _09573_ sky130_fd_sc_hd__nand2_1
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14244_ _06925_ _06932_ vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__nand2_1
XFILLER_32_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11456_ _03900_ _04164_ _04173_ _03954_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__o211a_1
XFILLER_109_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10407_ rbzero.tex_r1\[23\] rbzero.tex_r1\[24\] _03411_ vssd1 vssd1 vccd1 vccd1 _03416_
+ sky130_fd_sc_hd__mux2_1
X_14175_ _06435_ _06542_ _06847_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__o21ai_1
X_11387_ gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__clkbuf_4
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13126_ _05802_ _05813_ _05814_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__o21a_1
XFILLER_152_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10338_ _03379_ vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__clkbuf_1
X_18983_ rbzero.pov.spi_buffer\[39\] rbzero.pov.ready_buffer\[39\] _02651_ vssd1 vssd1
+ vccd1 vccd1 _02652_ sky130_fd_sc_hd__mux2_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _01500_ _01609_ _01714_ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__o21bai_2
XFILLER_152_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13057_ _05618_ _05745_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__and2_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10269_ rbzero.tex_b1\[24\] rbzero.tex_b1\[25\] _03333_ vssd1 vssd1 vccd1 vccd1 _03343_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12008_ net3 vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__buf_2
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17865_ _01646_ _01647_ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__xor2_2
XFILLER_120_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19604_ _07494_ _02955_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__nand2_1
XFILLER_66_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16816_ _09303_ _09358_ _09359_ _09282_ vssd1 vssd1 vccd1 vccd1 _09360_ sky130_fd_sc_hd__a31o_1
X_17796_ _01578_ _01579_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__xor2_1
XFILLER_226_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19535_ _02936_ vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13959_ _06646_ _06647_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__xnor2_1
X_16747_ _09296_ _09297_ _09295_ vssd1 vssd1 vccd1 vccd1 _09299_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16678_ rbzero.row_render.texu\[2\] _09260_ _09258_ rbzero.wall_tracer.texu\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__a22o_1
X_19466_ _02900_ vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__clkbuf_1
XFILLER_222_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18417_ rbzero.wall_tracer.rayAddendX\[-4\] _00013_ _02165_ _02169_ vssd1 vssd1 vccd1
+ vccd1 _00591_ sky130_fd_sc_hd__o22a_1
X_15629_ _08156_ _08242_ vssd1 vssd1 vccd1 vccd1 _08243_ sky130_fd_sc_hd__nor2_1
XFILLER_146_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19397_ _02863_ vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__clkinv_2
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18348_ _02101_ _02103_ _02102_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__o21ba_1
XFILLER_194_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18279_ _02048_ _02049_ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20310_ rbzero.traced_texVinit\[1\] _09266_ _08571_ _09261_ vssd1 vssd1 vccd1 vccd1
+ _01395_ sky130_fd_sc_hd__a22o_1
X_21290_ net133 _01306_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-12\] sky130_fd_sc_hd__dfxtp_1
Xinput50 i_tex_in[3] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_2
XFILLER_238_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20241_ _03253_ vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__clkinv_2
XFILLER_190_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20172_ _03197_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__inv_2
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11310_ _03784_ _03290_ _03293_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__o21a_1
X_20508_ net132 _00524_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-3\] sky130_fd_sc_hd__dfxtp_1
X_12290_ _04956_ _04957_ _04949_ _04983_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__or4_1
XFILLER_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11241_ rbzero.tex_r0\[45\] rbzero.tex_r0\[44\] _03959_ vssd1 vssd1 vccd1 vccd1 _03960_
+ sky130_fd_sc_hd__mux2_1
XTAP_7001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20439_ net138 _00470_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_7012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11172_ _03888_ _03890_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__nand2_1
XTAP_7056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15980_ _07388_ _08592_ _08067_ _07790_ vssd1 vssd1 vccd1 vccd1 _08593_ sky130_fd_sc_hd__or4_1
XTAP_6355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14931_ rbzero.wall_tracer.visualWallDist\[-2\] _07544_ _07408_ vssd1 vssd1 vccd1
+ vccd1 _07545_ sky130_fd_sc_hd__mux2_1
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17650_ _09833_ _07914_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__nor2_1
XFILLER_208_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14862_ _07426_ _07475_ vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__or2b_1
XFILLER_180_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16601_ _07680_ _08923_ vssd1 vssd1 vccd1 vccd1 _09210_ sky130_fd_sc_hd__nor2_1
X_13813_ _06499_ _06501_ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__or2b_1
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17581_ _10110_ _10116_ _10117_ vssd1 vssd1 vccd1 vccd1 _10118_ sky130_fd_sc_hd__nand3_1
XFILLER_180_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14793_ _07406_ rbzero.debug_overlay.playerY\[-4\] _05113_ vssd1 vssd1 vccd1 vccd1
+ _07407_ sky130_fd_sc_hd__mux2_1
XFILLER_17_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16532_ _08997_ _09000_ _08999_ vssd1 vssd1 vccd1 vccd1 _09141_ sky130_fd_sc_hd__a21bo_1
X_19320_ _02851_ vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13744_ _06420_ _06429_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__nor2_1
XFILLER_186_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10956_ rbzero.tex_b0\[21\] rbzero.tex_b0\[20\] _03704_ vssd1 vssd1 vccd1 vccd1 _03706_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16463_ _08937_ _08939_ vssd1 vssd1 vccd1 vccd1 _09073_ sky130_fd_sc_hd__nand2_1
XFILLER_204_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19251_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.new_leak\[4\] _02804_
+ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__mux2_1
XFILLER_108_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13675_ _06361_ _06363_ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__and2b_1
XFILLER_189_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10887_ _03669_ vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__clkbuf_1
XFILLER_231_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18202_ _01889_ _01891_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__nor2_1
X_15414_ _07981_ _07999_ _08001_ vssd1 vssd1 vccd1 vccd1 _08028_ sky130_fd_sc_hd__and3_1
XFILLER_148_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12626_ _05280_ _05286_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__nor2_1
X_19182_ _02768_ vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__clkbuf_1
XPHY_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16394_ _08869_ _08864_ vssd1 vssd1 vccd1 vccd1 _09004_ sky130_fd_sc_hd__and2b_1
XFILLER_188_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18133_ _01834_ _01913_ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__and2b_1
X_15345_ _07955_ _07957_ _07958_ vssd1 vssd1 vccd1 vccd1 _07959_ sky130_fd_sc_hd__a21o_1
XFILLER_223_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12557_ _05245_ _05150_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__nor2_1
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18064_ _01744_ _01844_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__xnor2_1
X_11508_ _04224_ _04225_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__nor2_1
X_15276_ _07552_ vssd1 vssd1 vccd1 vccd1 _07890_ sky130_fd_sc_hd__buf_2
X_12488_ _05168_ _05171_ _05173_ _05176_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__o211a_1
X_17015_ _09546_ _09555_ vssd1 vssd1 vccd1 vccd1 _09556_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14227_ _06101_ _06172_ _06542_ _06470_ vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__o22a_1
X_11439_ _03956_ _04139_ _04147_ _04156_ _03985_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__o311a_1
XFILLER_172_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14158_ _06642_ _06846_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13109_ _05795_ _05797_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__nor2_1
XFILLER_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14089_ _06754_ _06776_ _06777_ vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__a21bo_1
X_18966_ rbzero.pov.spi_buffer\[31\] rbzero.pov.ready_buffer\[31\] _02640_ vssd1 vssd1
+ vccd1 vccd1 _02643_ sky130_fd_sc_hd__mux2_1
XFILLER_79_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17917_ _01698_ _01699_ vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__and2_1
XFILLER_112_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18897_ rbzero.spi_registers.spi_counter\[6\] _02602_ _02605_ vssd1 vssd1 vccd1 vccd1
+ _00635_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17848_ _09428_ _08634_ _09463_ _08594_ vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__o22ai_1
XFILLER_82_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17779_ _01527_ _01562_ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__xor2_1
XFILLER_78_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19518_ _02927_ vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20790_ net102 _00806_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_vshift
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_241_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19449_ _02891_ vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__clkbuf_1
XFILLER_222_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21342_ _00365_ _01358_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21273_ _00322_ _01289_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20224_ rbzero.traced_texa\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _03241_
+ sky130_fd_sc_hd__nand2_1
XFILLER_11_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20155_ rbzero.traced_texa\[-2\] rbzero.texV\[-2\] vssd1 vssd1 vccd1 vccd1 _03183_
+ sky130_fd_sc_hd__and2_1
XFILLER_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20086_ _03131_ vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__clkinv_2
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _03629_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _04323_ _04502_ _04503_ _04504_ _03921_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__o221a_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20988_ net65 _01004_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10741_ _03592_ vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13460_ _06064_ _06060_ _06095_ _06066_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__a211o_1
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10672_ rbzero.tex_g1\[27\] rbzero.tex_g1\[28\] _03552_ vssd1 vssd1 vccd1 vccd1 _03557_
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12411_ _05059_ _05061_ _05103_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__nand3_1
XFILLER_220_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13391_ _06075_ _06079_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__xnor2_1
XFILLER_103_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15130_ _07442_ _07379_ _07400_ _07355_ vssd1 vssd1 vccd1 vccd1 _07744_ sky130_fd_sc_hd__o22ai_1
XFILLER_167_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12342_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__and2_1
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15061_ rbzero.wall_tracer.visualWallDist\[-10\] _03794_ vssd1 vssd1 vccd1 vccd1
+ _07675_ sky130_fd_sc_hd__nand2_2
XFILLER_142_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12273_ _04966_ rbzero.wall_tracer.trackDistY\[-10\] vssd1 vssd1 vccd1 vccd1 _04967_
+ sky130_fd_sc_hd__or2_1
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14012_ _06649_ _06700_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11224_ rbzero.tex_r0\[59\] _03939_ _03941_ _03942_ vssd1 vssd1 vccd1 vccd1 _03943_
+ sky130_fd_sc_hd__a31o_1
XFILLER_88_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18820_ _02523_ _02534_ _02539_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__nand3_1
XTAP_6130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11155_ rbzero.traced_texVinit\[8\] rbzero.spi_registers.vshift\[5\] vssd1 vssd1
+ vccd1 vccd1 _03874_ sky130_fd_sc_hd__nor2_1
XTAP_6141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18751_ _02443_ _02455_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__nand2_1
XTAP_6185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15963_ rbzero.debug_overlay.playerY\[-9\] rbzero.debug_overlay.playerX\[-9\] _07342_
+ vssd1 vssd1 vccd1 vccd1 _08577_ sky130_fd_sc_hd__mux2_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11086_ rbzero.wall_tracer.state\[14\] _03808_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__nand2_4
XFILLER_216_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17702_ _01485_ _01486_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__xor2_1
XTAP_5473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14914_ _07336_ _07527_ rbzero.wall_tracer.state\[13\] vssd1 vssd1 vccd1 vccd1 _07528_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_114_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15894_ _07424_ _08067_ _07520_ _08507_ vssd1 vssd1 vccd1 vccd1 _08508_ sky130_fd_sc_hd__a2bb2o_1
XTAP_5484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18682_ _02409_ _02410_ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__xor2_1
XTAP_5495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17633_ _10167_ _10168_ vssd1 vssd1 vccd1 vccd1 _10169_ sky130_fd_sc_hd__xnor2_1
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14845_ _07458_ rbzero.debug_overlay.playerY\[-7\] _05113_ vssd1 vssd1 vccd1 vccd1
+ _07459_ sky130_fd_sc_hd__mux2_1
XFILLER_223_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17564_ _08241_ _09463_ _09962_ _10100_ _09961_ vssd1 vssd1 vccd1 vccd1 _10101_ sky130_fd_sc_hd__o32a_1
X_14776_ _07389_ _07358_ vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__xnor2_1
XFILLER_223_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11988_ net15 net16 vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__and2b_1
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19303_ rbzero.pov.spi_counter\[0\] _02837_ _02838_ vssd1 vssd1 vccd1 vccd1 _02839_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_232_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16515_ _07878_ _08723_ vssd1 vssd1 vccd1 vccd1 _09124_ sky130_fd_sc_hd__nor2_1
X_13727_ _06408_ _06409_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__or2b_1
X_10939_ rbzero.tex_b0\[29\] rbzero.tex_b0\[28\] _03693_ vssd1 vssd1 vccd1 vccd1 _03697_
+ sky130_fd_sc_hd__mux2_1
XFILLER_205_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17495_ _09895_ _09897_ _09896_ vssd1 vssd1 vccd1 vccd1 _10032_ sky130_fd_sc_hd__o21ba_1
XFILLER_232_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19234_ _02799_ vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16446_ _07835_ _07680_ _08785_ _09055_ vssd1 vssd1 vccd1 vccd1 _09056_ sky130_fd_sc_hd__or4b_1
X_13658_ _06333_ _06340_ _06344_ _06346_ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__a22oi_1
XFILLER_231_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12609_ _05193_ _05297_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__xnor2_2
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16377_ _07792_ _07880_ _08717_ _08984_ vssd1 vssd1 vccd1 vccd1 _08987_ sky130_fd_sc_hd__or4_1
XFILLER_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19165_ rbzero.color_sky\[2\] _02752_ _02757_ vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__a21o_1
X_13589_ _06267_ _06276_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__and2_1
XFILLER_118_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18116_ _01774_ _01777_ _01895_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__nand3_1
X_15328_ _07762_ _07934_ _07941_ vssd1 vssd1 vccd1 vccd1 _07942_ sky130_fd_sc_hd__nand3_1
XFILLER_219_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19096_ rbzero.spi_registers.ss_buffer\[1\] rbzero.spi_registers.ss_buffer\[0\] _04920_
+ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__mux2_1
XFILLER_121_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18047_ _01827_ _01828_ _09275_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__o21a_1
X_15259_ _07869_ _07870_ _07872_ vssd1 vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__nand3_1
XFILLER_173_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19998_ _03122_ vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__clkinv_2
XFILLER_98_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18949_ rbzero.pov.spi_buffer\[23\] rbzero.pov.ready_buffer\[23\] _02629_ vssd1 vssd1
+ vccd1 vccd1 _02634_ sky130_fd_sc_hd__mux2_1
XFILLER_228_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20911_ net78 _00927_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_215_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20842_ _00060_ _00858_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20773_ net87 _00789_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout58 net59 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_2
XFILLER_167_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout69 net72 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21325_ _00348_ _01341_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21256_ _00305_ _01272_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20207_ rbzero.traced_texa\[6\] rbzero.texV\[6\] vssd1 vssd1 vccd1 vccd1 _03227_
+ sky130_fd_sc_hd__nand2_1
XFILLER_85_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21187_ _00236_ _01203_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_77_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20138_ _03163_ _03165_ _03164_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__o21bai_1
XFILLER_213_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ _05644_ _05648_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__xnor2_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20069_ _03129_ vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__clkinv_2
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11911_ net14 _04614_ _04617_ _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__and4b_1
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12891_ _05298_ _05300_ _05430_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__mux2_1
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ rbzero.wall_tracer.visualWallDist\[0\] _07252_ vssd1 vssd1 vccd1 vccd1 _07283_
+ sky130_fd_sc_hd__or2_1
XFILLER_2_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11842_ _04554_ _04555_ _03928_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__mux2_1
XFILLER_73_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _07230_ vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__clkbuf_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11773_ _04323_ _04485_ _04486_ _04487_ _03921_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__o221a_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _08786_ _08790_ _08909_ vssd1 vssd1 vccd1 vccd1 _08911_ sky130_fd_sc_hd__nand3_1
XFILLER_214_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13512_ _05553_ _05701_ _06200_ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__and3_1
XFILLER_53_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17280_ _09678_ _09689_ _09687_ vssd1 vssd1 vccd1 vccd1 _09819_ sky130_fd_sc_hd__a21oi_1
XFILLER_159_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ rbzero.tex_g1\[2\] rbzero.tex_g1\[3\] _03574_ vssd1 vssd1 vccd1 vccd1 _03584_
+ sky130_fd_sc_hd__mux2_1
XFILLER_213_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14492_ _05527_ _07141_ _07142_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__and3_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16231_ _08745_ _08713_ vssd1 vssd1 vccd1 vccd1 _08842_ sky130_fd_sc_hd__or2b_1
XFILLER_224_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13443_ _06122_ _05671_ _06028_ _05641_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10655_ rbzero.tex_g1\[35\] rbzero.tex_g1\[36\] _03541_ vssd1 vssd1 vccd1 vccd1 _03548_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16162_ _08618_ _08772_ _08773_ vssd1 vssd1 vccd1 vccd1 _08774_ sky130_fd_sc_hd__o21a_1
XFILLER_16_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13374_ _06061_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__or2b_1
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10586_ _03511_ vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__clkbuf_1
X_15113_ _07698_ _07661_ _07662_ _07726_ _07697_ vssd1 vssd1 vccd1 vccd1 _07727_ sky130_fd_sc_hd__a32o_1
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12325_ rbzero.wall_tracer.trackDistX\[-11\] _05018_ _04970_ vssd1 vssd1 vccd1 vccd1
+ _05019_ sky130_fd_sc_hd__o21ai_1
XFILLER_103_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16093_ _08704_ _08705_ vssd1 vssd1 vccd1 vccd1 _08706_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15044_ _07655_ _07657_ vssd1 vssd1 vccd1 vccd1 _07658_ sky130_fd_sc_hd__xnor2_2
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19921_ _03115_ vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__clkinv_2
XFILLER_177_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12256_ rbzero.wall_tracer.trackDistX\[-2\] vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__inv_2
XFILLER_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11207_ rbzero.tex_r0\[63\] rbzero.tex_r0\[62\] _03925_ vssd1 vssd1 vccd1 vccd1 _03926_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19852_ _03108_ vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__clkinv_2
X_12187_ _04883_ _04118_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__nor2_1
XFILLER_214_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18803_ _02522_ _02523_ vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__nand2_1
XFILLER_150_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11138_ rbzero.traced_texVinit\[2\] rbzero.texV\[2\] rbzero.texV\[1\] rbzero.traced_texVinit\[1\]
+ _03856_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__a221o_1
XFILLER_96_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19783_ _04628_ _03813_ _02717_ _03085_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__a22o_1
XFILLER_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16995_ _08890_ _08718_ _08985_ _08596_ vssd1 vssd1 vccd1 vccd1 _09536_ sky130_fd_sc_hd__o22ai_1
XFILLER_49_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18734_ _02443_ _02446_ _02457_ _09256_ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a31o_1
X_15946_ _08557_ _08559_ vssd1 vssd1 vccd1 vccd1 _08560_ sky130_fd_sc_hd__xor2_1
XTAP_5270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11069_ rbzero.wall_tracer.state\[13\] vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__clkinv_2
XTAP_5281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18665_ rbzero.wall_tracer.rayAddendY\[-4\] _00013_ _02392_ _02395_ vssd1 vssd1 vccd1
+ vccd1 _00613_ sky130_fd_sc_hd__o22a_1
XFILLER_237_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15877_ _08488_ _08489_ _08490_ vssd1 vssd1 vccd1 vccd1 _08491_ sky130_fd_sc_hd__nand3_1
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17616_ _09903_ _09905_ _10046_ _10044_ vssd1 vssd1 vccd1 vccd1 _10152_ sky130_fd_sc_hd__a31o_1
XFILLER_188_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14828_ _07439_ _07440_ _07441_ vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__a21o_1
XFILLER_184_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18596_ _02275_ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__inv_2
XFILLER_221_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17547_ _10080_ _10082_ vssd1 vssd1 vccd1 vccd1 _10084_ sky130_fd_sc_hd__and2_1
X_14759_ _07372_ _05203_ _05210_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__and3b_1
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17478_ _09881_ _09776_ vssd1 vssd1 vccd1 vccd1 _10016_ sky130_fd_sc_hd__or2b_1
XFILLER_220_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19217_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.new_sky\[3\] _02786_
+ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__mux2_1
X_16429_ _08771_ _08636_ vssd1 vssd1 vccd1 vccd1 _09039_ sky130_fd_sc_hd__nand2_1
XFILLER_242_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19148_ rbzero.floor_leak\[1\] _02744_ _02747_ _02738_ vssd1 vssd1 vccd1 vccd1 _00744_
+ sky130_fd_sc_hd__o211a_1
XFILLER_160_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19079_ _02589_ _02576_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__nand2_1
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21110_ _00159_ _01126_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21041_ _00090_ _01057_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20825_ _00043_ _00841_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_243_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20756_ net106 _00772_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20687_ net76 _00703_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[67\] sky130_fd_sc_hd__dfxtp_1
XFILLER_206_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10440_ _03388_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__clkbuf_4
XFILLER_104_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10371_ rbzero.tex_r1\[40\] rbzero.tex_r1\[41\] _03389_ vssd1 vssd1 vccd1 vccd1 _03397_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12110_ _04797_ _04808_ _04817_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__a21o_1
X_21308_ net114 _01324_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13090_ _05762_ _05778_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__xor2_1
XFILLER_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12041_ net3 net4 vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__nor2_1
X_21239_ _00288_ _01255_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15800_ _08377_ _08385_ _08382_ vssd1 vssd1 vccd1 vccd1 _08414_ sky130_fd_sc_hd__a21o_1
XFILLER_63_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13992_ _06633_ _06680_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__xnor2_1
X_16780_ _09325_ _09326_ _09327_ vssd1 vssd1 vccd1 vccd1 _09328_ sky130_fd_sc_hd__or3_1
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15731_ _08330_ _08344_ vssd1 vssd1 vccd1 vccd1 _08345_ sky130_fd_sc_hd__nor2_1
X_12943_ _05624_ _05631_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__nor2_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ _02198_ _02199_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__nand2_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _08274_ _07971_ _08275_ vssd1 vssd1 vccd1 vccd1 _08276_ sky130_fd_sc_hd__o21a_1
X_12874_ _05559_ _05562_ _05480_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _09937_ _09938_ vssd1 vssd1 vccd1 vccd1 _09939_ sky130_fd_sc_hd__xor2_1
XFILLER_185_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ rbzero.wall_tracer.trackDistX\[-5\] rbzero.wall_tracer.trackDistY\[-5\] _07258_
+ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__mux2_1
X_11825_ _03909_ _04536_ _04537_ _04538_ _03920_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__o221a_1
X_18381_ rbzero.wall_tracer.trackDistY\[11\] rbzero.wall_tracer.stepDistY\[11\] vssd1
+ vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__xor2_1
X_15593_ _08198_ _08205_ vssd1 vssd1 vccd1 vccd1 _08207_ sky130_fd_sc_hd__nor2_1
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17332_ _09740_ _09742_ vssd1 vssd1 vccd1 vccd1 _09871_ sky130_fd_sc_hd__or2b_1
X_14544_ _07213_ _07216_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__nand2_1
XFILLER_159_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _03968_ _04468_ _04469_ _04470_ _03972_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__o221a_1
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10707_ _03575_ vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__clkbuf_1
X_17263_ _09800_ _09801_ vssd1 vssd1 vccd1 vccd1 _09802_ sky130_fd_sc_hd__xor2_1
XFILLER_202_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14475_ _05527_ _07113_ _05577_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__a21o_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11687_ rbzero.tex_g1\[9\] rbzero.tex_g1\[8\] _03980_ vssd1 vssd1 vccd1 vccd1 _04403_
+ sky130_fd_sc_hd__mux2_1
X_19002_ _02661_ vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16214_ _08711_ _08824_ vssd1 vssd1 vccd1 vccd1 _08826_ sky130_fd_sc_hd__or2_1
X_13426_ _05618_ _05745_ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__nand2_2
XFILLER_31_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17194_ _09474_ vssd1 vssd1 vccd1 vccd1 _09734_ sky130_fd_sc_hd__inv_2
X_10638_ rbzero.tex_g1\[43\] rbzero.tex_g1\[44\] _03530_ vssd1 vssd1 vccd1 vccd1 _03539_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16145_ _08755_ _08756_ vssd1 vssd1 vccd1 vccd1 _08757_ sky130_fd_sc_hd__nand2_1
XFILLER_31_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13357_ _06044_ _06045_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10569_ rbzero.tex_r0\[13\] rbzero.tex_r0\[12\] _03501_ vssd1 vssd1 vccd1 vccd1 _03503_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12308_ rbzero.wall_tracer.trackDistY\[5\] vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__inv_2
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16076_ _08686_ _08688_ vssd1 vssd1 vccd1 vccd1 _08689_ sky130_fd_sc_hd__or2_1
XFILLER_143_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13288_ _05948_ _05975_ _05976_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__a21boi_1
X_15027_ _07466_ rbzero.wall_tracer.stepDistX\[1\] vssd1 vssd1 vccd1 vccd1 _07641_
+ sky130_fd_sc_hd__nand2_1
X_19904_ _03113_ vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__clkinv_2
XFILLER_170_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12239_ _04933_ _03730_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__nor2_1
XFILLER_64_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19835_ _03106_ vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__clkinv_2
XFILLER_69_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19766_ _04246_ _04628_ _04631_ _03074_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__or4_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16978_ _09387_ _09390_ _09518_ vssd1 vssd1 vccd1 vccd1 _09519_ sky130_fd_sc_hd__o21a_1
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput4 i_gpout0_sel[1] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_4
XFILLER_237_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18717_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__nand2_1
X_15929_ _08541_ _08542_ vssd1 vssd1 vccd1 vccd1 _08543_ sky130_fd_sc_hd__nand2_1
XFILLER_83_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19697_ rbzero.debug_overlay.playerY\[4\] _02834_ _03043_ rbzero.debug_overlay.playerY\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__or4b_1
XFILLER_36_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18648_ _02373_ _02378_ _02379_ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__o21ai_1
XFILLER_188_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18579_ _02275_ rbzero.wall_tracer.rayAddendX\[8\] vssd1 vssd1 vccd1 vccd1 _02320_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_149_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20610_ net92 _00626_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_221_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20541_ net137 _00557_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20472_ net111 _00488_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21024_ net109 _01040_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11610_ _04323_ _04324_ _04325_ _04326_ _03923_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__o221a_1
XFILLER_58_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20808_ _00026_ _00824_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12590_ _03816_ _05069_ _05112_ _05278_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__a31o_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11541_ rbzero.debug_overlay.vplaneX\[10\] _04236_ _04258_ vssd1 vssd1 vccd1 vccd1
+ _04259_ sky130_fd_sc_hd__a21o_1
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20739_ net107 _00755_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14260_ _06844_ _06935_ _06946_ _06948_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__a31o_1
XFILLER_183_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11472_ _03924_ _04185_ _04189_ _03899_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__a211o_1
XFILLER_184_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13211_ _05890_ _05891_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__nand2_1
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10423_ _03424_ vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__clkbuf_1
X_14191_ _06843_ _06876_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__nand2_1
XFILLER_125_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13142_ _05815_ _05816_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__nor2_1
XFILLER_152_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10354_ _03387_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_191_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17950_ _01730_ _01731_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__or2_1
X_13073_ _05724_ _05732_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__nand2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10285_ _03351_ vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16901_ _09426_ _09194_ _09442_ vssd1 vssd1 vccd1 vccd1 _09443_ sky130_fd_sc_hd__a21o_1
X_12024_ _03294_ _03295_ gpout0.vpos\[8\] _04110_ net3 _04731_ vssd1 vssd1 vccd1 vccd1
+ _04733_ sky130_fd_sc_hd__mux4_1
XFILLER_26_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17881_ _01661_ _01662_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__nand2_1
XFILLER_61_1318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19620_ rbzero.pov.ready_buffer\[70\] _02963_ _02981_ _02992_ vssd1 vssd1 vccd1 vccd1
+ _02993_ sky130_fd_sc_hd__o211a_1
XFILLER_78_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16832_ _09124_ _09125_ vssd1 vssd1 vccd1 vccd1 _09374_ sky130_fd_sc_hd__nand2_1
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19551_ _02944_ vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16763_ _09304_ _09306_ _09305_ vssd1 vssd1 vccd1 vccd1 _09313_ sky130_fd_sc_hd__a21boi_1
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13975_ _06663_ _06645_ vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18502_ _02247_ rbzero.wall_tracer.rayAddendX\[3\] vssd1 vssd1 vccd1 vccd1 _02248_
+ sky130_fd_sc_hd__nand2_1
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15714_ _08325_ _08327_ vssd1 vssd1 vccd1 vccd1 _08328_ sky130_fd_sc_hd__or2b_1
XFILLER_206_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12926_ _05613_ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__nor2_2
X_19482_ _02908_ vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16694_ _09254_ vssd1 vssd1 vccd1 vccd1 _09264_ sky130_fd_sc_hd__buf_2
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18433_ _02172_ _02176_ _02173_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__o21ai_1
XFILLER_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15645_ _08255_ _08257_ _08258_ vssd1 vssd1 vccd1 vccd1 _08259_ sky130_fd_sc_hd__a21oi_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12857_ _05537_ _05545_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__nor2_1
XFILLER_146_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18364_ _02121_ _02122_ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11808_ _04520_ _04521_ _03908_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__mux2_1
XFILLER_221_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12788_ _05459_ _05445_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__and2_1
X_15576_ _08179_ _08185_ _08187_ vssd1 vssd1 vccd1 vccd1 _08190_ sky130_fd_sc_hd__and3_1
XFILLER_159_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _09852_ _09853_ vssd1 vssd1 vccd1 vccd1 _09854_ sky130_fd_sc_hd__xnor2_1
XFILLER_226_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14527_ _07203_ vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11739_ _04323_ _04451_ _04452_ _04453_ _03972_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__o221a_1
X_18295_ rbzero.wall_tracer.trackDistY\[-2\] _02039_ _02063_ _09354_ vssd1 vssd1 vccd1
+ vccd1 _00575_ sky130_fd_sc_hd__o22a_1
XFILLER_222_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17246_ _09777_ _09778_ _09784_ vssd1 vssd1 vccd1 vccd1 _09785_ sky130_fd_sc_hd__a21oi_1
XFILLER_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14458_ _05577_ _07143_ _07144_ _07133_ vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__o31ai_1
XFILLER_128_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13409_ _06087_ _06097_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__and2_1
X_17177_ _09698_ _09716_ vssd1 vssd1 vccd1 vccd1 _09717_ sky130_fd_sc_hd__xor2_1
X_14389_ _06990_ _07045_ _07077_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__a21oi_1
XFILLER_183_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16128_ _08667_ _08679_ _08677_ vssd1 vssd1 vccd1 vccd1 _08740_ sky130_fd_sc_hd__a21oi_1
XFILLER_196_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16059_ _07880_ _07621_ _08671_ _07792_ vssd1 vssd1 vccd1 vccd1 _08672_ sky130_fd_sc_hd__o22ai_1
XFILLER_142_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19818_ _03105_ vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__clkinv_2
XFILLER_233_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19749_ rbzero.pov.ready_buffer\[21\] _03069_ _03070_ _02275_ _02832_ vssd1 vssd1
+ vccd1 vccd1 _01022_ sky130_fd_sc_hd__o221a_1
XFILLER_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_20 rbzero.traced_texa\[-11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_31 net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_42 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20524_ net96 _00540_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.wall\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20455_ net97 _00016_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20386_ net131 _00417_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21007_ net79 _01023_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_88_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13760_ _06430_ _06448_ _06446_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10972_ rbzero.tex_b0\[13\] rbzero.tex_b0\[12\] _03704_ vssd1 vssd1 vccd1 vccd1 _03714_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12711_ _05336_ _05361_ _05363_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__or3_1
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13691_ _06376_ _06379_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__nor2_1
XFILLER_95_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15430_ _08043_ _07966_ vssd1 vssd1 vccd1 vccd1 _08044_ sky130_fd_sc_hd__xnor2_1
X_12642_ _05295_ _05330_ _05271_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__and3_1
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15361_ _07468_ _07388_ _07973_ _07974_ vssd1 vssd1 vccd1 vccd1 _07975_ sky130_fd_sc_hd__o31a_1
X_12573_ rbzero.wall_tracer.rcp_sel\[0\] _05242_ _05244_ _05249_ _05261_ vssd1 vssd1
+ vccd1 vccd1 _05262_ sky130_fd_sc_hd__a2111o_1
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17100_ _07332_ _09640_ vssd1 vssd1 vccd1 vccd1 _09641_ sky130_fd_sc_hd__and2_1
XFILLER_50_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14312_ _06999_ _07000_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11524_ _04208_ _04241_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__nor2_2
X_18080_ _01859_ _01860_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__xor2_1
XFILLER_200_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15292_ _07782_ _07813_ _07904_ _07905_ vssd1 vssd1 vccd1 vccd1 _07906_ sky130_fd_sc_hd__o211ai_1
XFILLER_7_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17031_ _08595_ _09571_ _07817_ _08594_ vssd1 vssd1 vccd1 vccd1 _09572_ sky130_fd_sc_hd__o22ai_1
X_14243_ _06923_ _06924_ vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__or2_1
XFILLER_172_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11455_ _03972_ _04167_ _04172_ _03950_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__a211o_1
XFILLER_194_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10406_ _03415_ vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__clkbuf_1
X_14174_ _06101_ _06423_ _06858_ _06862_ vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__o31a_1
XFILLER_152_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11386_ _04104_ _04101_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__nand2_1
XFILLER_152_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13125_ _05786_ _05801_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__nand2_1
XFILLER_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10337_ rbzero.tex_r1\[56\] rbzero.tex_r1\[57\] _03377_ vssd1 vssd1 vccd1 vccd1 _03379_
+ sky130_fd_sc_hd__mux2_1
X_18982_ _02607_ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__clkbuf_4
XFILLER_124_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17933_ _10023_ _10024_ _01501_ _01715_ vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__a31o_2
X_13056_ _05526_ _05546_ _05553_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a21o_2
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ _03342_ vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12007_ o_rgb[6] _04669_ _04685_ _04716_ vssd1 vssd1 vccd1 vccd1 o_gpout[2] sky130_fd_sc_hd__o22a_2
XFILLER_239_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17864_ _01583_ _01594_ _01593_ vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__a21oi_2
XFILLER_230_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10199_ _03306_ vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19603_ rbzero.pov.ready_buffer\[67\] _07564_ _02962_ vssd1 vssd1 vccd1 vccd1 _02979_
+ sky130_fd_sc_hd__mux2_1
XFILLER_226_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16815_ _09355_ _09356_ _09357_ vssd1 vssd1 vccd1 vccd1 _09359_ sky130_fd_sc_hd__o21ai_1
XFILLER_238_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17795_ _09968_ _09197_ _01459_ _01461_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__o31a_1
XFILLER_66_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19534_ rbzero.pov.spi_buffer\[62\] rbzero.pov.spi_buffer\[63\] _02932_ vssd1 vssd1
+ vccd1 vccd1 _02936_ sky130_fd_sc_hd__mux2_1
XFILLER_207_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16746_ _09295_ _09296_ _09297_ vssd1 vssd1 vccd1 vccd1 _09298_ sky130_fd_sc_hd__or3_1
X_13958_ _06595_ _06597_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__xor2_1
XFILLER_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12909_ _05406_ _05530_ _05597_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__o21ai_1
X_19465_ rbzero.pov.spi_buffer\[29\] rbzero.pov.spi_buffer\[30\] _02899_ vssd1 vssd1
+ vccd1 vccd1 _02900_ sky130_fd_sc_hd__mux2_1
XFILLER_222_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16677_ rbzero.row_render.texu\[1\] _09260_ _09258_ rbzero.wall_tracer.texu\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__a22o_1
X_13889_ _05767_ _06483_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__or2_1
XFILLER_59_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18416_ _02166_ _02167_ _02168_ _09254_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a31o_1
X_15628_ _08240_ _07986_ _08060_ _08241_ vssd1 vssd1 vccd1 vccd1 _08242_ sky130_fd_sc_hd__o22a_1
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19396_ _02863_ vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__clkinv_2
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18347_ rbzero.wall_tracer.trackDistY\[6\] rbzero.wall_tracer.stepDistY\[6\] vssd1
+ vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__and2_1
XFILLER_194_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15559_ _08161_ _08164_ vssd1 vssd1 vccd1 vccd1 _08173_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18278_ _02040_ _02042_ _02041_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__a21boi_1
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput40 i_mode[1] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_8
X_17229_ _09766_ _09767_ _09768_ vssd1 vssd1 vccd1 vccd1 _09769_ sky130_fd_sc_hd__and3_1
XFILLER_174_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput51 i_vec_csb vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_4
XFILLER_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20240_ _03253_ vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__clkinv_2
XFILLER_192_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20171_ _03193_ _03194_ _03195_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__and3_1
XFILLER_131_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20507_ net132 _00523_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11240_ _03925_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__clkbuf_4
X_20438_ net139 _00469_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11171_ _03880_ _03889_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20369_ net92 _00402_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.c6 sky130_fd_sc_hd__dfxtp_2
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14930_ _07543_ rbzero.debug_overlay.playerY\[-2\] _05113_ vssd1 vssd1 vccd1 vccd1
+ _07544_ sky130_fd_sc_hd__mux2_1
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14861_ _07456_ _07474_ vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__nand2_1
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16600_ _09114_ _09208_ vssd1 vssd1 vccd1 vccd1 _09209_ sky130_fd_sc_hd__xnor2_1
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ _06491_ _06493_ _06500_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__o21ai_1
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17580_ _10114_ _10115_ _10111_ vssd1 vssd1 vccd1 vccd1 _10117_ sky130_fd_sc_hd__a21o_1
XFILLER_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14792_ _07404_ _07405_ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__and2_1
XFILLER_235_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16531_ _09138_ _09139_ vssd1 vssd1 vccd1 vccd1 _09140_ sky130_fd_sc_hd__and2_1
XFILLER_217_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13743_ _06395_ _06431_ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__or2_1
X_10955_ _03705_ vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19250_ _02808_ vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__clkbuf_1
X_16462_ _09069_ _09070_ _09046_ vssd1 vssd1 vccd1 vccd1 _09072_ sky130_fd_sc_hd__a21o_1
XFILLER_189_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13674_ _06316_ _06362_ _06323_ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__o21ba_1
XFILLER_32_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10886_ rbzero.tex_b0\[54\] rbzero.tex_b0\[53\] _03660_ vssd1 vssd1 vccd1 vccd1 _03669_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18201_ _01974_ _01980_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15413_ _08004_ _08026_ vssd1 vssd1 vccd1 vccd1 _08027_ sky130_fd_sc_hd__xor2_1
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ _05281_ _05313_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__xnor2_2
X_19181_ _09247_ _02767_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__and2_1
XPHY_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16393_ _08995_ _09002_ vssd1 vssd1 vccd1 vccd1 _09003_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18132_ _01911_ _01912_ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__or2_1
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15344_ _07931_ _07954_ vssd1 vssd1 vccd1 vccd1 _07958_ sky130_fd_sc_hd__nor2_1
XFILLER_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12556_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__and2_1
XFILLER_156_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11507_ _04199_ _04220_ _04196_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__or3b_2
X_18063_ _09968_ _09976_ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__nor2_1
XFILLER_156_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15275_ _07355_ _07387_ _07552_ _07550_ vssd1 vssd1 vccd1 vccd1 _07889_ sky130_fd_sc_hd__or4_1
XFILLER_184_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12487_ _05174_ _05175_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__and2_1
XFILLER_32_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17014_ _09553_ _09554_ vssd1 vssd1 vccd1 vccd1 _09555_ sky130_fd_sc_hd__and2b_1
X_14226_ _05959_ _06483_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__nor2_1
X_11438_ _03921_ _04151_ _04155_ _03898_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__a211o_1
XFILLER_137_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14157_ _05740_ _06483_ vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__nor2_1
XFILLER_140_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11369_ rbzero.row_render.size\[1\] _04086_ _04087_ _04042_ vssd1 vssd1 vccd1 vccd1
+ _04088_ sky130_fd_sc_hd__a31o_1
XFILLER_119_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13108_ _05673_ _05796_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__xor2_1
X_14088_ _06755_ _06756_ _06775_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__nand3_1
XFILLER_119_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18965_ _02642_ vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__clkbuf_1
XFILLER_239_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17916_ _01691_ _01692_ _01697_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__nand3_1
X_13039_ _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__clkbuf_2
XFILLER_26_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18896_ rbzero.spi_registers.spi_counter\[6\] _02602_ _02589_ vssd1 vssd1 vccd1 vccd1
+ _02605_ sky130_fd_sc_hd__o21ai_1
XTAP_6890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17847_ _08594_ _09428_ _08634_ _09462_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__or4_1
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17778_ _01547_ _01561_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19517_ rbzero.pov.spi_buffer\[54\] rbzero.pov.spi_buffer\[55\] _02921_ vssd1 vssd1
+ vccd1 vccd1 _02927_ sky130_fd_sc_hd__mux2_1
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16729_ _09282_ vssd1 vssd1 vccd1 vccd1 _09283_ sky130_fd_sc_hd__clkbuf_4
XFILLER_35_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19448_ rbzero.pov.spi_buffer\[21\] rbzero.pov.spi_buffer\[22\] _02888_ vssd1 vssd1
+ vccd1 vccd1 _02891_ sky130_fd_sc_hd__mux2_1
XFILLER_126_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19379_ _02860_ vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__clkinv_2
XFILLER_206_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21341_ _00364_ _01357_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21272_ _00321_ _01288_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20223_ rbzero.traced_texa\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _03240_
+ sky130_fd_sc_hd__or2_1
XFILLER_78_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20154_ rbzero.traced_texa\[-2\] rbzero.texV\[-2\] vssd1 vssd1 vccd1 vccd1 _03182_
+ sky130_fd_sc_hd__nor2_1
XFILLER_131_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20085_ _03131_ vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__clkinv_2
XFILLER_131_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20987_ net65 _01003_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10740_ rbzero.tex_g0\[59\] rbzero.tex_g0\[58\] _03512_ vssd1 vssd1 vccd1 vccd1 _03592_
+ sky130_fd_sc_hd__mux2_1
XFILLER_129_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10671_ _03556_ vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ _05056_ _05058_ _05063_ _05064_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__a211o_1
XFILLER_51_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13390_ _06042_ _06076_ _06077_ _06078_ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__o22ai_2
XFILLER_138_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12341_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__nor2_1
XFILLER_142_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15060_ _07672_ _07673_ _07646_ vssd1 vssd1 vccd1 vccd1 _07674_ sky130_fd_sc_hd__a21o_1
X_12272_ rbzero.wall_tracer.trackDistX\[-10\] vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__inv_2
XFILLER_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14011_ _06313_ _06483_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__nor2_1
XFILLER_181_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11223_ _03915_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__buf_4
XFILLER_135_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11154_ rbzero.traced_texVinit\[8\] rbzero.spi_registers.vshift\[5\] vssd1 vssd1
+ vccd1 vccd1 _03873_ sky130_fd_sc_hd__and2_1
XFILLER_175_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18750_ _02472_ rbzero.wall_tracer.rayAddendY\[3\] vssd1 vssd1 vccd1 vccd1 _02474_
+ sky130_fd_sc_hd__or2_1
XTAP_6175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15962_ _08454_ _08456_ vssd1 vssd1 vccd1 vccd1 _08576_ sky130_fd_sc_hd__xor2_2
X_11085_ _03802_ _03807_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__nor2_4
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17701_ _10109_ _10127_ _10126_ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__a21boi_1
XTAP_6197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14913_ rbzero.wall_tracer.rayAddendY\[-3\] rbzero.wall_tracer.rayAddendX\[-3\] rbzero.wall_tracer.side
+ vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__mux2_1
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18681_ _02398_ _02402_ _02399_ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__o21ai_1
X_15893_ _08296_ vssd1 vssd1 vccd1 vccd1 _08507_ sky130_fd_sc_hd__clkinv_2
XTAP_5485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17632_ _08750_ _09114_ vssd1 vssd1 vccd1 vccd1 _10168_ sky130_fd_sc_hd__nor2_1
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14844_ _07357_ _07457_ vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__and2_1
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17563_ _08787_ _09207_ _08240_ vssd1 vssd1 vccd1 vccd1 _10100_ sky130_fd_sc_hd__a21oi_1
XFILLER_217_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14775_ rbzero.debug_overlay.playerY\[-5\] vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__inv_2
X_11987_ net16 net15 vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__and2b_1
XFILLER_186_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19302_ rbzero.pov.ss_buffer\[1\] _03442_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__nor2_2
XFILLER_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16514_ _09033_ _09015_ vssd1 vssd1 vccd1 vccd1 _09123_ sky130_fd_sc_hd__or2b_1
XFILLER_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13726_ _06326_ _06411_ _06414_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__a21boi_1
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17494_ rbzero.wall_tracer.trackDistX\[5\] rbzero.wall_tracer.stepDistX\[5\] vssd1
+ vssd1 vccd1 vccd1 _10031_ sky130_fd_sc_hd__and2_1
X_10938_ _03696_ vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__clkbuf_1
XFILLER_220_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19233_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.new_floor\[3\]
+ _02795_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__mux2_1
X_16445_ rbzero.wall_tracer.stepDistX\[7\] _08633_ _04929_ vssd1 vssd1 vccd1 vccd1
+ _09055_ sky130_fd_sc_hd__mux2_4
XFILLER_189_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13657_ _06333_ _06340_ _06345_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__a21oi_2
X_10869_ _03604_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__clkbuf_4
XFILLER_158_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12608_ _05277_ _05289_ _05292_ _05296_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__o31a_1
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19164_ rbzero.spi_registers.new_sky\[2\] rbzero.spi_registers.got_new_sky _02724_
+ _02753_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__a31o_1
XFILLER_223_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16376_ _07880_ _08717_ _08985_ _07878_ vssd1 vssd1 vccd1 vccd1 _08986_ sky130_fd_sc_hd__o22a_1
XFILLER_160_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13588_ _06267_ _06276_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__nor2_1
X_18115_ _01774_ _01777_ _01895_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a21o_1
XFILLER_118_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15327_ _07938_ _07939_ _07940_ vssd1 vssd1 vccd1 vccd1 _07941_ sky130_fd_sc_hd__a21bo_1
XFILLER_158_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12539_ rbzero.wall_tracer.visualWallDist\[-4\] _05189_ rbzero.wall_tracer.rcp_sel\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__a21o_1
XFILLER_145_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19095_ _02711_ vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18046_ _01824_ _01825_ _01826_ _09351_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__a31o_1
XFILLER_117_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15258_ _07741_ _07755_ _07871_ vssd1 vssd1 vccd1 vccd1 _07872_ sky130_fd_sc_hd__a21o_1
XFILLER_172_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14209_ _06887_ _06897_ vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__or2b_1
X_15189_ _07485_ _07567_ vssd1 vssd1 vccd1 vccd1 _07803_ sky130_fd_sc_hd__or2_1
XFILLER_141_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19997_ _03122_ vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__clkinv_2
XFILLER_141_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18948_ _02633_ vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18879_ _02590_ _02591_ _02592_ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__and3_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20910_ net61 _00926_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20841_ _00059_ _00857_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20772_ net103 _00788_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_leak
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_223_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout59 net73 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21324_ _00347_ _01340_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21255_ _00304_ _01271_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20206_ rbzero.traced_texa\[6\] rbzero.texV\[6\] vssd1 vssd1 vccd1 vccd1 _03226_
+ sky130_fd_sc_hd__nor2_1
XFILLER_132_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21186_ _00235_ _01202_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20137_ rbzero.traced_texa\[-5\] rbzero.texV\[-5\] vssd1 vssd1 vccd1 vccd1 _03168_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_137_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20068_ _03129_ vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__clkinv_2
XFILLER_218_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _04618_ net11 _04620_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__and3_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12890_ _05517_ _05578_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__nand2_1
XFILLER_73_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11841_ rbzero.tex_b1\[17\] rbzero.tex_b1\[16\] _04544_ vssd1 vssd1 vccd1 vccd1 _04555_
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14560_ rbzero.wall_tracer.stepDistY\[7\] _07229_ _04925_ vssd1 vssd1 vccd1 vccd1
+ _07230_ sky130_fd_sc_hd__mux2_1
XFILLER_198_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11772_ rbzero.tex_b0\[31\] _04143_ _04145_ _03930_ vssd1 vssd1 vccd1 vccd1 _04487_
+ sky130_fd_sc_hd__a31o_1
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13511_ _06198_ _06199_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _03583_ vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14491_ _07133_ _07007_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__nor2_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _08664_ _08727_ vssd1 vssd1 vccd1 vccd1 _08841_ sky130_fd_sc_hd__or2b_1
XFILLER_220_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13442_ _06028_ _05612_ _05625_ _05715_ _06130_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__a41o_1
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10654_ _03547_ vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16161_ _08046_ _07837_ _08617_ vssd1 vssd1 vccd1 vccd1 _08773_ sky130_fd_sc_hd__a21o_1
X_13373_ _06027_ _06059_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__xor2_1
XFILLER_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10585_ rbzero.tex_r0\[5\] rbzero.tex_r0\[4\] _03501_ vssd1 vssd1 vccd1 vccd1 _03511_
+ sky130_fd_sc_hd__mux2_1
XFILLER_177_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15112_ _07709_ _07710_ vssd1 vssd1 vccd1 vccd1 _07726_ sky130_fd_sc_hd__nand2_1
X_12324_ rbzero.wall_tracer.trackDistY\[-11\] vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__inv_2
XFILLER_186_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16092_ _08567_ _08582_ _08565_ vssd1 vssd1 vccd1 vccd1 _08705_ sky130_fd_sc_hd__o21a_1
XFILLER_170_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15043_ _07446_ _07448_ _07656_ _07447_ vssd1 vssd1 vccd1 vccd1 _07657_ sky130_fd_sc_hd__o211a_1
X_12255_ _04947_ rbzero.wall_tracer.trackDistY\[-3\] rbzero.wall_tracer.trackDistY\[-4\]
+ _04948_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__a22o_1
XFILLER_154_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19920_ _03115_ vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__clkinv_2
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11206_ _03903_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__buf_4
XFILLER_68_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19851_ _03108_ vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__clkinv_2
XFILLER_69_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12186_ net37 _04890_ _04891_ net36 vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__a31o_1
XFILLER_123_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11137_ rbzero.traced_texVinit\[1\] rbzero.texV\[1\] rbzero.texV\[0\] rbzero.traced_texVinit\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__o211a_1
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18802_ _04260_ _02498_ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__nand2_1
X_19782_ _03073_ _03086_ _03087_ vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16994_ _09533_ _09534_ vssd1 vssd1 vccd1 vccd1 _09535_ sky130_fd_sc_hd__and2_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18733_ _02443_ _02446_ _02457_ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__a21oi_1
X_15945_ _07640_ _07960_ _08558_ vssd1 vssd1 vccd1 vccd1 _08559_ sky130_fd_sc_hd__a21oi_1
XTAP_5260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11068_ _03790_ _03791_ _03792_ _03730_ rbzero.wall_tracer.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _00011_ sky130_fd_sc_hd__a311o_1
XFILLER_114_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18664_ _02166_ _02393_ _02394_ _09254_ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__a31o_1
XFILLER_236_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15876_ _07839_ _07844_ _07836_ vssd1 vssd1 vccd1 vccd1 _08490_ sky130_fd_sc_hd__a21bo_1
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17615_ _10141_ _10038_ vssd1 vssd1 vccd1 vccd1 _10151_ sky130_fd_sc_hd__or2b_1
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14827_ _04927_ rbzero.wall_tracer.stepDistX\[-3\] vssd1 vssd1 vccd1 vccd1 _07441_
+ sky130_fd_sc_hd__nor2_1
XFILLER_188_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18595_ rbzero.wall_tracer.rayAddendX\[9\] _03812_ _09269_ _02332_ _02334_ vssd1
+ vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__o221a_1
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17546_ _10080_ _10082_ vssd1 vssd1 vccd1 vccd1 _10083_ sky130_fd_sc_hd__nor2_1
XFILLER_205_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14758_ _07371_ _05267_ _05215_ vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__or3b_1
XFILLER_205_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13709_ _06383_ _06397_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__and2_1
XFILLER_177_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17477_ _09900_ _10014_ vssd1 vssd1 vccd1 vccd1 _10015_ sky130_fd_sc_hd__xor2_1
X_14689_ rbzero.wall_tracer.stepDistX\[-1\] _07199_ _07316_ vssd1 vssd1 vccd1 vccd1
+ _07319_ sky130_fd_sc_hd__mux2_1
XFILLER_225_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19216_ _02789_ vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__clkbuf_1
X_16428_ _07696_ _08640_ _08272_ vssd1 vssd1 vccd1 vccd1 _09038_ sky130_fd_sc_hd__a21o_1
XFILLER_220_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19147_ rbzero.spi_registers.new_leak\[1\] _02745_ vssd1 vssd1 vccd1 vccd1 _02747_
+ sky130_fd_sc_hd__or2_1
X_16359_ _08880_ _08847_ vssd1 vssd1 vccd1 vccd1 _08969_ sky130_fd_sc_hd__or2b_1
XFILLER_146_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19078_ _02701_ vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18029_ _01695_ _01810_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__xor2_1
X_21040_ _00089_ _01056_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20824_ _00042_ _00840_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20755_ net106 _00771_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20686_ net76 _00702_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[66\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10370_ _03396_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21307_ net133 _01323_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12040_ net3 _04718_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__and2_1
XFILLER_46_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21238_ _00287_ _01254_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21169_ _00218_ _01185_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13991_ _06658_ _06678_ _06679_ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__a21oi_1
XFILLER_150_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15730_ _08289_ _08329_ _08328_ _08324_ vssd1 vssd1 vccd1 vccd1 _08344_ sky130_fd_sc_hd__o211a_1
XFILLER_111_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12942_ _05626_ _05630_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__and2_1
XFILLER_86_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15661_ _07435_ _07507_ vssd1 vssd1 vccd1 vccd1 _08275_ sky130_fd_sc_hd__or2_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12873_ _05501_ _05529_ _05561_ _05405_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__o211a_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _09429_ _07914_ vssd1 vssd1 vccd1 vccd1 _09938_ sky130_fd_sc_hd__nor2_1
XFILLER_2_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _07245_ _07269_ _07270_ _07251_ vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__o211a_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ rbzero.wall_tracer.trackDistY\[10\] rbzero.wall_tracer.stepDistY\[10\] _02133_
+ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__a21o_1
X_11824_ rbzero.tex_b1\[47\] _03938_ _03940_ _03915_ vssd1 vssd1 vccd1 vccd1 _04538_
+ sky130_fd_sc_hd__a31o_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _08198_ _08205_ vssd1 vssd1 vccd1 vccd1 _08206_ sky130_fd_sc_hd__xor2_2
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _09848_ _09869_ vssd1 vssd1 vccd1 vccd1 _09870_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _07174_ _07092_ _07215_ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__a21oi_1
XFILLER_159_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ rbzero.tex_b0\[41\] _04143_ _04145_ _03957_ vssd1 vssd1 vccd1 vccd1 _04470_
+ sky130_fd_sc_hd__a31o_1
XFILLER_222_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17262_ _08890_ _08725_ vssd1 vssd1 vccd1 vccd1 _09801_ sky130_fd_sc_hd__nor2_1
XFILLER_109_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10706_ rbzero.tex_g1\[11\] rbzero.tex_g1\[12\] _03574_ vssd1 vssd1 vccd1 vccd1 _03575_
+ sky130_fd_sc_hd__mux2_1
X_14474_ _05602_ _05408_ vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__nand2_1
X_11686_ _04400_ _04401_ _03997_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__mux2_1
XFILLER_202_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19001_ rbzero.pov.spi_buffer\[48\] rbzero.pov.ready_buffer\[48\] _02651_ vssd1 vssd1
+ vccd1 vccd1 _02661_ sky130_fd_sc_hd__mux2_1
X_16213_ _08711_ _08824_ vssd1 vssd1 vccd1 vccd1 _08825_ sky130_fd_sc_hd__nand2_1
XFILLER_122_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13425_ _06099_ _06100_ _06113_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__and3_1
X_17193_ _09474_ _09476_ _09609_ _09732_ vssd1 vssd1 vccd1 vccd1 _09733_ sky130_fd_sc_hd__or4bb_2
XFILLER_128_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10637_ _03538_ vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16144_ _08240_ _07712_ _07736_ _08241_ vssd1 vssd1 vccd1 vccd1 _08756_ sky130_fd_sc_hd__o22ai_1
XFILLER_128_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13356_ _05537_ _05627_ _05657_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__or3_1
X_10568_ _03502_ vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12307_ rbzero.wall_tracer.trackDistY\[4\] vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__inv_2
X_16075_ _08529_ _08552_ _08687_ vssd1 vssd1 vccd1 vccd1 _08688_ sky130_fd_sc_hd__a21oi_1
X_13287_ _05974_ _05950_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__or2b_1
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10499_ rbzero.tex_r0\[46\] rbzero.tex_r0\[45\] _03457_ vssd1 vssd1 vccd1 vccd1 _03466_
+ sky130_fd_sc_hd__mux2_1
XFILLER_216_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15026_ _07588_ _07615_ _07639_ vssd1 vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__a21oi_2
X_19903_ _02862_ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__buf_4
XFILLER_190_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12238_ _04932_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__clkbuf_8
XFILLER_155_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12169_ net34 net35 net36 vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__a21o_1
X_19834_ _03106_ vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__clkinv_2
XFILLER_233_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16977_ _09385_ _09386_ vssd1 vssd1 vccd1 vccd1 _09518_ sky130_fd_sc_hd__nand2_1
X_19765_ _04110_ _04106_ _03073_ _04114_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__or4_1
XFILLER_81_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 i_gpout0_sel[2] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_4
X_15928_ _07881_ _07885_ _08540_ vssd1 vssd1 vccd1 vccd1 _08542_ sky130_fd_sc_hd__nand3_1
XFILLER_42_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18716_ _02428_ rbzero.wall_tracer.rayAddendY\[0\] vssd1 vssd1 vccd1 vccd1 _02442_
+ sky130_fd_sc_hd__or2_1
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19696_ _03048_ _03051_ _03003_ vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__a21oi_1
XFILLER_237_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18647_ rbzero.debug_overlay.vplaneY\[-7\] rbzero.wall_tracer.rayAddendY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__nand2_1
X_15859_ _07453_ rbzero.wall_tracer.stepDistY\[6\] vssd1 vssd1 vccd1 vccd1 _08473_
+ sky130_fd_sc_hd__nand2_1
XFILLER_225_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18578_ _02308_ _02312_ _02317_ _03818_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__a31o_1
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17529_ _10062_ _10064_ vssd1 vssd1 vccd1 vccd1 _10066_ sky130_fd_sc_hd__nand2_1
XFILLER_127_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20540_ net123 _00556_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20471_ net111 _00487_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21023_ net110 _01039_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20807_ _00025_ _00823_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_243_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11540_ rbzero.debug_overlay.vplaneX\[-9\] _04240_ _04253_ _04257_ vssd1 vssd1 vccd1
+ vccd1 _04258_ sky130_fd_sc_hd__a211o_1
XFILLER_106_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20738_ net105 _00754_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ _04186_ _04187_ _04188_ _03957_ _03946_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__o221a_1
XFILLER_168_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20669_ net74 _00685_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13210_ _05715_ _05749_ _05893_ _05898_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__o31a_1
XFILLER_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10422_ rbzero.tex_r1\[16\] rbzero.tex_r1\[17\] _03422_ vssd1 vssd1 vccd1 vccd1 _03424_
+ sky130_fd_sc_hd__mux2_1
X_14190_ _06839_ _06835_ _06838_ _06878_ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__a211oi_1
XFILLER_104_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13141_ _05825_ _05829_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__xor2_1
X_10353_ rbzero.tex_r1\[48\] rbzero.tex_r1\[49\] _03377_ vssd1 vssd1 vccd1 vccd1 _03387_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13072_ _05758_ _05760_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10284_ rbzero.tex_b1\[17\] rbzero.tex_b1\[18\] _03344_ vssd1 vssd1 vccd1 vccd1 _03351_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16900_ _09433_ _09441_ vssd1 vssd1 vccd1 vccd1 _09442_ sky130_fd_sc_hd__xnor2_1
XFILLER_215_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12023_ gpout0.hpos\[2\] _04080_ _04628_ _04101_ net3 _04731_ vssd1 vssd1 vccd1 vccd1
+ _04732_ sky130_fd_sc_hd__mux4_1
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17880_ _01661_ _01662_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__or2_1
XFILLER_238_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16831_ _08979_ vssd1 vssd1 vccd1 vccd1 _09373_ sky130_fd_sc_hd__clkbuf_4
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19550_ rbzero.pov.spi_buffer\[70\] rbzero.pov.spi_buffer\[71\] _02865_ vssd1 vssd1
+ vccd1 vccd1 _02944_ sky130_fd_sc_hd__mux2_1
XFILLER_232_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16762_ rbzero.wall_tracer.trackDistX\[-8\] rbzero.wall_tracer.stepDistX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _09312_ sky130_fd_sc_hd__and2_1
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13974_ _06407_ _06642_ _06644_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__a21bo_1
XFILLER_20_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18501_ rbzero.debug_overlay.vplaneX\[10\] vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__buf_2
XFILLER_207_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15713_ _08324_ _08326_ vssd1 vssd1 vccd1 vccd1 _08327_ sky130_fd_sc_hd__and2_1
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12925_ _05537_ _05545_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__or2_1
X_19481_ rbzero.pov.spi_buffer\[37\] rbzero.pov.spi_buffer\[38\] _02899_ vssd1 vssd1
+ vccd1 vccd1 _02908_ sky130_fd_sc_hd__mux2_1
XFILLER_74_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16693_ rbzero.traced_texa\[-3\] _09262_ _09263_ rbzero.wall_tracer.visualWallDist\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__a22o_1
XFILLER_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18432_ _02181_ _02182_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__nand2_1
XFILLER_98_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15644_ _08253_ _08254_ vssd1 vssd1 vccd1 vccd1 _08258_ sky130_fd_sc_hd__nor2_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _05538_ _05541_ _05544_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__o21a_2
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18363_ _02113_ _02115_ _02114_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__a21boi_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ rbzero.tex_b1\[51\] rbzero.tex_b1\[50\] _04032_ vssd1 vssd1 vccd1 vccd1 _04521_
+ sky130_fd_sc_hd__mux2_1
X_15575_ _08148_ _08158_ vssd1 vssd1 vccd1 vccd1 _08189_ sky130_fd_sc_hd__xnor2_2
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12787_ _05381_ _05395_ _05253_ _05378_ _05462_ _05463_ vssd1 vssd1 vccd1 vccd1 _05476_
+ sky130_fd_sc_hd__mux4_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _09182_ _09197_ vssd1 vssd1 vccd1 vccd1 _09853_ sky130_fd_sc_hd__nor2_1
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14526_ rbzero.wall_tracer.stepDistY\[0\] _07202_ _07193_ vssd1 vssd1 vccd1 vccd1
+ _07203_ sky130_fd_sc_hd__mux2_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18294_ _01997_ _02061_ _02062_ _02013_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__a31o_1
X_11738_ rbzero.tex_b0\[59\] _04143_ _04145_ _03930_ vssd1 vssd1 vccd1 vccd1 _04453_
+ sky130_fd_sc_hd__a31o_1
XFILLER_226_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17245_ _09782_ _09783_ vssd1 vssd1 vccd1 vccd1 _09784_ sky130_fd_sc_hd__nand2_1
X_14457_ _07115_ _07111_ _07114_ _07130_ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__a22o_1
XFILLER_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11669_ rbzero.tex_g1\[17\] rbzero.tex_g1\[16\] _04378_ vssd1 vssd1 vccd1 vccd1 _04385_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13408_ _06085_ _06086_ vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__or2_1
X_17176_ _09699_ _09715_ vssd1 vssd1 vccd1 vccd1 _09716_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14388_ _06987_ _07032_ _07033_ _07036_ _07029_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__o311a_1
XFILLER_116_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16127_ _08729_ _08738_ vssd1 vssd1 vccd1 vccd1 _08739_ sky130_fd_sc_hd__xnor2_1
XFILLER_192_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13339_ _05488_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__clkbuf_4
XFILLER_143_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16058_ _08670_ vssd1 vssd1 vccd1 vccd1 _08671_ sky130_fd_sc_hd__clkbuf_4
XFILLER_157_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15009_ _07616_ _07618_ _07622_ vssd1 vssd1 vccd1 vccd1 _07623_ sky130_fd_sc_hd__nor3_1
XFILLER_237_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19817_ _03105_ vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__clkinv_2
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19748_ rbzero.pov.ready_buffer\[20\] _03067_ _03068_ rbzero.debug_overlay.vplaneX\[0\]
+ _03015_ vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__a221o_1
XFILLER_84_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19679_ rbzero.pov.ready_buffer\[54\] _02963_ _03012_ _03037_ vssd1 vssd1 vccd1 vccd1
+ _03038_ sky130_fd_sc_hd__o211a_1
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_10 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 rbzero.wall_tracer.visualWallDist\[-3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_32 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20523_ net96 _00539_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.wall\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_43 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20454_ net118 _00005_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20385_ net131 _00416_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21006_ net82 _01022_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10971_ _03713_ vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12710_ _05360_ _05393_ _05397_ _05398_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__and4_1
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13690_ _06377_ _06378_ _06324_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__a21boi_1
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12641_ _05200_ _05201_ _05203_ _03790_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__a22o_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15360_ _07969_ _07972_ vssd1 vssd1 vccd1 vccd1 _07974_ sky130_fd_sc_hd__or2_1
XFILLER_157_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12572_ _05256_ _05260_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__or2_1
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14311_ _06690_ _06970_ _06971_ vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__a21boi_1
XFILLER_178_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11523_ _04078_ _04221_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__nand2_1
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15291_ _07873_ _07874_ _07903_ vssd1 vssd1 vccd1 vccd1 _07905_ sky130_fd_sc_hd__a21o_1
XFILLER_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17030_ _07672_ vssd1 vssd1 vccd1 vccd1 _09571_ sky130_fd_sc_hd__buf_2
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14242_ _06908_ _06927_ _06930_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__nand3_1
XFILLER_144_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11454_ _03957_ _04169_ _04170_ _04171_ _03923_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__o221a_1
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10405_ rbzero.tex_r1\[24\] rbzero.tex_r1\[25\] _03411_ vssd1 vssd1 vccd1 vccd1 _03415_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14173_ _05959_ _06389_ _06861_ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__or3b_1
X_11385_ gpout0.vpos\[5\] vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__buf_2
XFILLER_139_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13124_ _05808_ _05812_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10336_ _03378_ vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18981_ _02650_ vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__clkbuf_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17932_ _01502_ _01714_ vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__or2_1
X_13055_ _05653_ _05655_ _05642_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__a21bo_1
XFILLER_139_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ rbzero.tex_b1\[25\] rbzero.tex_b1\[26\] _03333_ vssd1 vssd1 vccd1 vccd1 _03342_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12006_ _04688_ _04690_ _04693_ _04715_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__a31o_1
X_17863_ _01625_ _01645_ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__xnor2_2
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10198_ rbzero.tex_b1\[58\] rbzero.tex_b1\[59\] _03300_ vssd1 vssd1 vccd1 vccd1 _03306_
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19602_ _02956_ _02976_ _02977_ _02978_ vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__o211a_1
XFILLER_213_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16814_ _09355_ _09356_ _09357_ vssd1 vssd1 vccd1 vccd1 _09358_ sky130_fd_sc_hd__or3_1
X_17794_ _01576_ _01577_ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__xor2_1
XFILLER_238_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16745_ rbzero.wall_tracer.trackDistX\[-10\] rbzero.wall_tracer.stepDistX\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _09297_ sky130_fd_sc_hd__and2_1
X_19533_ _02935_ vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__clkbuf_1
X_13957_ _06407_ _06642_ _06644_ _06645_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__a22o_1
XFILLER_34_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12908_ _05531_ _05586_ _05472_ _05569_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__o31ai_1
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19464_ _02865_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__clkbuf_4
XFILLER_234_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16676_ rbzero.row_render.texu\[0\] _09260_ _09258_ rbzero.wall_tracer.texu\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__a22o_1
XFILLER_234_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13888_ _06543_ _06544_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__xor2_1
XFILLER_34_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15627_ _07800_ vssd1 vssd1 vccd1 vccd1 _08241_ sky130_fd_sc_hd__buf_4
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18415_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__or2_1
XFILLER_222_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12839_ _05378_ _05381_ _05448_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__mux2_1
X_19395_ _02863_ vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__clkinv_2
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18346_ rbzero.wall_tracer.trackDistY\[6\] rbzero.wall_tracer.stepDistY\[6\] vssd1
+ vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__nor2_1
X_15558_ _08114_ _08166_ vssd1 vssd1 vccd1 vccd1 _08172_ sky130_fd_sc_hd__xnor2_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14509_ rbzero.wall_tracer.stepDistY\[-4\] _07189_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _07190_ sky130_fd_sc_hd__mux2_1
XFILLER_187_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18277_ _02046_ _02047_ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__and2b_1
XFILLER_148_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15489_ _08073_ _08102_ vssd1 vssd1 vccd1 vccd1 _08103_ sky130_fd_sc_hd__nor2_1
XFILLER_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17228_ _09643_ _09647_ vssd1 vssd1 vccd1 vccd1 _09768_ sky130_fd_sc_hd__nand2_1
Xinput30 i_gpout4_sel[3] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_6
Xinput41 i_mode[2] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_8
Xinput52 i_vec_mosi vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_8
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17159_ _09590_ _09600_ _09598_ vssd1 vssd1 vccd1 vccd1 _09699_ sky130_fd_sc_hd__a21oi_1
XFILLER_162_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20170_ _03193_ _03194_ _03195_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__a21o_1
XFILLER_107_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20506_ net132 _00522_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20437_ net135 _00468_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11170_ rbzero.traced_texVinit\[11\] rbzero.texV\[11\] vssd1 vssd1 vccd1 vccd1 _03889_
+ sky130_fd_sc_hd__xnor2_1
XTAP_7025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20368_ net92 _00401_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.d6 sky130_fd_sc_hd__dfxtp_2
XTAP_7036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20299_ _03258_ vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__clkinv_2
XTAP_6346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14860_ _07468_ _07469_ _07456_ _07473_ vssd1 vssd1 vccd1 vccd1 _07474_ sky130_fd_sc_hd__or4bb_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ _06489_ _06494_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__or2b_1
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14791_ rbzero.debug_overlay.playerY\[-5\] _07358_ rbzero.debug_overlay.playerY\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__o21ai_1
XFILLER_112_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16530_ _09128_ _09137_ vssd1 vssd1 vccd1 vccd1 _09139_ sky130_fd_sc_hd__or2_1
XFILLER_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13742_ _06374_ _06394_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__and2_1
XFILLER_147_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10954_ rbzero.tex_b0\[22\] rbzero.tex_b0\[21\] _03704_ vssd1 vssd1 vccd1 vccd1 _03705_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16461_ _09046_ _09069_ _09070_ vssd1 vssd1 vccd1 vccd1 _09071_ sky130_fd_sc_hd__nand3_1
X_13673_ _05722_ _06306_ _06318_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__o21a_1
XFILLER_147_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10885_ _03668_ vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__clkbuf_1
X_18200_ _01976_ _01979_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__xnor2_1
XFILLER_223_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15412_ _08023_ _08024_ _08025_ vssd1 vssd1 vccd1 vccd1 _08026_ sky130_fd_sc_hd__a21oi_1
XFILLER_227_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12624_ _05277_ _05312_ _05286_ _05305_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__o31ai_2
X_19180_ rbzero.spi_registers.new_floor\[2\] rbzero.color_floor\[2\] _02763_ vssd1
+ vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__mux2_1
XPHY_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16392_ _08996_ _09001_ vssd1 vssd1 vccd1 vccd1 _09002_ sky130_fd_sc_hd__xnor2_1
XPHY_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18131_ _01908_ _01910_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__and2_1
XFILLER_145_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15343_ _07640_ _07956_ vssd1 vssd1 vccd1 vccd1 _07957_ sky130_fd_sc_hd__nor2_1
XPHY_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12555_ _05189_ _05093_ _05243_ _05219_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__o211a_1
XFILLER_196_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18062_ _09968_ _09978_ _01744_ _01637_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__o31a_1
X_11506_ _03783_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__inv_2
XFILLER_117_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15274_ _07885_ _07887_ vssd1 vssd1 vccd1 vccd1 _07888_ sky130_fd_sc_hd__and2_1
X_12486_ rbzero.debug_overlay.facingX\[-1\] rbzero.wall_tracer.rayAddendX\[7\] vssd1
+ vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__or2_1
XFILLER_156_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17013_ _09547_ _09552_ vssd1 vssd1 vccd1 vccd1 _09554_ sky130_fd_sc_hd__or2_1
XFILLER_32_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14225_ _06470_ _06172_ vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__or2_1
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11437_ _03910_ _04152_ _04153_ _04154_ _03945_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__o221a_1
XFILLER_158_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14156_ _06643_ _06844_ vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__nand2_1
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11368_ gpout0.hpos\[1\] gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__or2_1
XFILLER_28_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13107_ _05627_ _05604_ _05657_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__or3_1
XFILLER_113_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10319_ _03369_ vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__clkbuf_1
X_14087_ _06755_ _06756_ _06775_ vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__a21o_1
XFILLER_193_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18964_ rbzero.pov.spi_buffer\[30\] rbzero.pov.ready_buffer\[30\] _02640_ vssd1 vssd1
+ vccd1 vccd1 _02642_ sky130_fd_sc_hd__mux2_1
XFILLER_234_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11299_ rbzero.tex_r0\[5\] rbzero.tex_r0\[4\] _03961_ vssd1 vssd1 vccd1 vccd1 _04018_
+ sky130_fd_sc_hd__mux2_1
XFILLER_224_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17915_ _01691_ _01692_ _01697_ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__a21o_1
X_13038_ _05703_ _05704_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__and2_1
XFILLER_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18895_ _02604_ vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__clkbuf_1
XTAP_6880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17846_ _01584_ _01588_ _01628_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__a21bo_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17777_ _01559_ _01560_ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__and2b_1
X_14989_ _07598_ _07602_ vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__nor2_1
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19516_ _02926_ vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__clkbuf_1
X_16728_ _05026_ _09272_ vssd1 vssd1 vccd1 vccd1 _09282_ sky130_fd_sc_hd__nand2_4
XFILLER_165_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19447_ _02890_ vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__clkbuf_1
X_16659_ _09256_ _03809_ vssd1 vssd1 vccd1 vccd1 _09257_ sky130_fd_sc_hd__nor2_8
XFILLER_165_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19378_ _02860_ vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__clkinv_2
XFILLER_72_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18329_ _02089_ _02090_ _02091_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__nand3_1
XFILLER_176_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21340_ _00363_ _01356_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21271_ _00320_ _01287_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20222_ rbzero.texV\[8\] _03137_ _03142_ _03239_ vssd1 vssd1 vccd1 vccd1 _01326_
+ sky130_fd_sc_hd__a22o_1
XFILLER_116_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20153_ _03093_ _03180_ _03181_ _03064_ rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1
+ _01315_ sky130_fd_sc_hd__a32o_1
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20084_ _03131_ vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__clkinv_2
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20986_ net65 _01002_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10670_ rbzero.tex_g1\[28\] rbzero.tex_g1\[29\] _03552_ vssd1 vssd1 vccd1 vccd1 _03556_
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12340_ _05031_ _05032_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__nand2_1
XFILLER_166_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12271_ rbzero.wall_tracer.trackDistX\[-9\] vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__inv_2
XFILLER_153_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ _06266_ _06542_ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__or2_1
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11222_ _03940_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__clkbuf_4
XFILLER_175_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11153_ _03840_ _03868_ _03871_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__o21a_1
XTAP_6121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15961_ _08574_ _07431_ _07343_ vssd1 vssd1 vccd1 vccd1 _08575_ sky130_fd_sc_hd__mux2_1
X_11084_ _03803_ _03290_ _03806_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__or3b_2
XTAP_6165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17700_ _01470_ _01484_ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__xnor2_1
XFILLER_216_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14912_ _07100_ _07135_ _07336_ vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__a21o_1
XTAP_5464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15892_ _07424_ _08296_ _07591_ _07790_ vssd1 vssd1 vccd1 vccd1 _08506_ sky130_fd_sc_hd__or4_1
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18680_ _02407_ _02408_ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__nand2_1
XTAP_5475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17631_ _10165_ _10166_ vssd1 vssd1 vccd1 vccd1 _10167_ sky130_fd_sc_hd__or2b_1
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerY\[-9\] rbzero.debug_overlay.playerY\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__o21ai_1
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17562_ _10097_ _10098_ vssd1 vssd1 vccd1 vccd1 _10099_ sky130_fd_sc_hd__xnor2_1
XFILLER_205_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14774_ _07387_ vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__buf_2
XFILLER_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11986_ gpout2.clk_div\[1\] _04667_ _04695_ _04115_ vssd1 vssd1 vccd1 vccd1 _04696_
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16513_ _09032_ _09016_ vssd1 vssd1 vccd1 vccd1 _09122_ sky130_fd_sc_hd__or2b_1
XFILLER_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19301_ rbzero.pov.sclk_buffer\[2\] rbzero.pov.sclk_buffer\[1\] vssd1 vssd1 vccd1
+ vccd1 _02837_ sky130_fd_sc_hd__nor2b_2
X_13725_ _06412_ _06413_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__or2b_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17493_ rbzero.wall_tracer.trackDistX\[5\] rbzero.wall_tracer.stepDistX\[5\] vssd1
+ vssd1 vccd1 vccd1 _10030_ sky130_fd_sc_hd__nor2_1
XFILLER_182_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10937_ rbzero.tex_b0\[30\] rbzero.tex_b0\[29\] _03693_ vssd1 vssd1 vccd1 vccd1 _03696_
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16444_ _09047_ _09053_ vssd1 vssd1 vccd1 vccd1 _09054_ sky130_fd_sc_hd__xnor2_1
XFILLER_220_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19232_ _02798_ vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13656_ _05818_ _06321_ _06331_ _06317_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_182_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10868_ _03659_ vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12607_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__buf_2
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19163_ _02756_ vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__clkbuf_1
X_16375_ _08984_ vssd1 vssd1 vccd1 vccd1 _08985_ sky130_fd_sc_hd__buf_2
XFILLER_157_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13587_ _06242_ _06275_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__xnor2_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10799_ _03623_ vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18114_ _08123_ _09115_ _01764_ _01762_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__o31a_1
XFILLER_160_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15326_ _07936_ _07718_ _07935_ vssd1 vssd1 vccd1 vccd1 _07940_ sky130_fd_sc_hd__or3_1
XFILLER_158_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12538_ _05219_ _05226_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__or2_1
X_19094_ net42 rbzero.spi_registers.ss_buffer\[0\] _02708_ vssd1 vssd1 vccd1 vccd1
+ _02711_ sky130_fd_sc_hd__mux2_1
XFILLER_157_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18045_ _01824_ _01825_ _01826_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__a21oi_1
X_15257_ _07715_ _07740_ vssd1 vssd1 vccd1 vccd1 _07871_ sky130_fd_sc_hd__nor2_1
XFILLER_172_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12469_ _05156_ _05157_ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__nand2_2
X_14208_ _06862_ _06888_ _06892_ _06894_ _06896_ vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__a32o_1
XFILLER_126_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15188_ _07799_ _07801_ vssd1 vssd1 vccd1 vccd1 _07802_ sky130_fd_sc_hd__nand2_1
XFILLER_119_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14139_ _06827_ _06806_ vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__xor2_1
XFILLER_119_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19996_ _03122_ vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__clkinv_2
XFILLER_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18947_ rbzero.pov.spi_buffer\[22\] rbzero.pov.ready_buffer\[22\] _02629_ vssd1 vssd1
+ vccd1 vccd1 _02633_ sky130_fd_sc_hd__mux2_1
XFILLER_98_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18878_ rbzero.spi_registers.spi_counter\[0\] _02576_ rbzero.spi_registers.spi_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__a21o_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17829_ rbzero.wall_tracer.trackDistX\[7\] rbzero.wall_tracer.stepDistX\[7\] vssd1
+ vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__or2_1
XFILLER_227_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20840_ _00058_ _00856_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20771_ net103 _00787_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21323_ _00346_ _01339_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21254_ _00303_ _01270_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20205_ rbzero.texV\[5\] _03137_ _03142_ _03225_ vssd1 vssd1 vccd1 vccd1 _01323_
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21185_ _00234_ _01201_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20136_ _03093_ _03166_ _03167_ _03137_ rbzero.texV\[-6\] vssd1 vssd1 vccd1 vccd1
+ _01312_ sky130_fd_sc_hd__a32o_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20067_ _03129_ vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__clkinv_2
XFILLER_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ rbzero.tex_b1\[19\] rbzero.tex_b1\[18\] _04544_ vssd1 vssd1 vccd1 vccd1 _04554_
+ sky130_fd_sc_hd__mux2_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11771_ rbzero.tex_b0\[30\] _03962_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__and2_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20969_ net71 _00985_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13510_ _05608_ _05767_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__nor2_1
XFILLER_159_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ rbzero.tex_g1\[3\] rbzero.tex_g1\[4\] _03574_ vssd1 vssd1 vccd1 vccd1 _03583_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14490_ _07173_ vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__clkbuf_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13441_ _05629_ _06129_ _06109_ _06108_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__o211a_1
XFILLER_55_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10653_ rbzero.tex_g1\[36\] rbzero.tex_g1\[37\] _03541_ vssd1 vssd1 vccd1 vccd1 _03547_
+ sky130_fd_sc_hd__mux2_1
XFILLER_224_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16160_ _08771_ _07837_ vssd1 vssd1 vccd1 vccd1 _08772_ sky130_fd_sc_hd__nand2_1
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13372_ _06029_ _06036_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__or2_1
XFILLER_194_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10584_ _03510_ vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15111_ _07470_ _07443_ _07663_ _07711_ vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__or4_1
XFILLER_186_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12323_ _05016_ rbzero.wall_tracer.trackDistX\[-8\] _04976_ _04978_ vssd1 vssd1 vccd1
+ vccd1 _05017_ sky130_fd_sc_hd__a211o_1
XFILLER_103_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16091_ _08702_ _08703_ vssd1 vssd1 vccd1 vccd1 _08704_ sky130_fd_sc_hd__or2_1
XFILLER_182_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15042_ _07028_ _07076_ _07098_ _07133_ vssd1 vssd1 vccd1 vccd1 _07656_ sky130_fd_sc_hd__a31o_1
XFILLER_142_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12254_ rbzero.wall_tracer.trackDistX\[-4\] vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__inv_2
XFILLER_155_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11205_ _03923_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__buf_4
XFILLER_194_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19850_ _03108_ vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__clkinv_2
XFILLER_64_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12185_ _04883_ _04447_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__nand2_1
X_18801_ _02520_ _02521_ _02498_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__a21o_1
XFILLER_205_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11136_ rbzero.texV\[3\] _03854_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__xor2_1
XFILLER_150_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19781_ _04632_ _04631_ _03808_ _02753_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__a31o_1
X_16993_ _09531_ _09532_ vssd1 vssd1 vccd1 vccd1 _09534_ sky130_fd_sc_hd__or2_1
XFILLER_27_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18732_ _02455_ _02456_ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__nand2_1
XFILLER_209_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15944_ _07928_ _07929_ _07959_ vssd1 vssd1 vccd1 vccd1 _08558_ sky130_fd_sc_hd__and3_1
XTAP_5250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11067_ rbzero.wall_tracer.state\[11\] vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__inv_2
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15875_ _07827_ _07847_ _08486_ _08487_ vssd1 vssd1 vccd1 vccd1 _08489_ sky130_fd_sc_hd__a2bb2o_1
XTAP_5294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18663_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__nand2_1
XFILLER_97_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17614_ _10139_ _10140_ vssd1 vssd1 vccd1 vccd1 _10150_ sky130_fd_sc_hd__or2_1
XFILLER_221_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14826_ rbzero.wall_tracer.state\[13\] rbzero.wall_tracer.stepDistY\[-3\] rbzero.wall_tracer.state\[6\]
+ vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__a21oi_2
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18594_ _02315_ _02318_ _02333_ _03818_ vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__a211o_1
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17545_ _09933_ _09940_ _10081_ vssd1 vssd1 vccd1 vccd1 _10082_ sky130_fd_sc_hd__a21oi_1
X_14757_ _05226_ _07370_ _05221_ _05230_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__or4b_1
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11969_ _04677_ _04678_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__or2_1
XFILLER_189_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13708_ _06395_ _06396_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__xor2_1
X_17476_ _10011_ _10013_ vssd1 vssd1 vccd1 vccd1 _10014_ sky130_fd_sc_hd__xnor2_1
XFILLER_162_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14688_ _07318_ vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19215_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.new_sky\[2\] _02786_
+ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__mux2_1
X_16427_ _08046_ _08636_ vssd1 vssd1 vccd1 vccd1 _09037_ sky130_fd_sc_hd__and2_1
X_13639_ _06309_ _06327_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__or2_1
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16358_ _08838_ _08962_ _08967_ vssd1 vssd1 vccd1 vccd1 _08968_ sky130_fd_sc_hd__a21o_1
XFILLER_121_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19146_ rbzero.floor_leak\[0\] _02744_ _02746_ _02738_ vssd1 vssd1 vccd1 vccd1 _00743_
+ sky130_fd_sc_hd__o211a_1
XFILLER_203_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15309_ _07921_ _07922_ vssd1 vssd1 vccd1 vccd1 _07923_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16289_ _08898_ _08899_ vssd1 vssd1 vccd1 vccd1 _08900_ sky130_fd_sc_hd__xor2_2
XFILLER_12_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19077_ rbzero.spi_registers.spi_buffer\[10\] rbzero.spi_registers.spi_buffer\[9\]
+ _02689_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__mux2_1
XFILLER_146_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18028_ _01808_ _01809_ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__nor2_1
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19979_ _03120_ vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__clkinv_2
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20823_ _00041_ _00839_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20754_ net106 _00770_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20685_ net76 _00701_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[65\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21306_ net132 _01322_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_174_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21237_ _00286_ _01253_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21168_ _00217_ _01184_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20119_ rbzero.traced_texa\[-8\] rbzero.texV\[-8\] vssd1 vssd1 vccd1 vccd1 _03153_
+ sky130_fd_sc_hd__nor2_1
X_13990_ _06659_ _06677_ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__nor2_1
X_21099_ _00148_ _01115_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_246_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12941_ _05627_ _05629_ _05525_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__or3_2
XFILLER_46_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15660_ _08202_ vssd1 vssd1 vccd1 vccd1 _08274_ sky130_fd_sc_hd__clkbuf_4
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _05501_ _05560_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__nand2_1
XFILLER_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14611_ rbzero.wall_tracer.visualWallDist\[-6\] _07249_ vssd1 vssd1 vccd1 vccd1 _07270_
+ sky130_fd_sc_hd__or2_1
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ rbzero.tex_b1\[46\] _04119_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__and2_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _08201_ _08203_ _08204_ vssd1 vssd1 vccd1 vccd1 _08205_ sky130_fd_sc_hd__a21oi_2
XFILLER_2_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17330_ _09866_ _09868_ vssd1 vssd1 vccd1 vccd1 _09869_ sky130_fd_sc_hd__xor2_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14542_ _07075_ _07088_ _07214_ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ rbzero.tex_b0\[40\] _03962_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__and2_1
XFILLER_186_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _09798_ _09799_ vssd1 vssd1 vccd1 vccd1 _09800_ sky130_fd_sc_hd__or2b_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _03298_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__clkbuf_4
XFILLER_202_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14473_ _07158_ vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11685_ rbzero.tex_g1\[13\] rbzero.tex_g1\[12\] _03980_ vssd1 vssd1 vccd1 vccd1 _04401_
+ sky130_fd_sc_hd__mux2_1
XFILLER_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16212_ _08822_ _08823_ vssd1 vssd1 vccd1 vccd1 _08824_ sky130_fd_sc_hd__xor2_1
X_19000_ _02660_ vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__clkbuf_1
X_13424_ _06104_ _06105_ _06111_ _06112_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__a31o_1
XFILLER_146_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17192_ _04939_ _09200_ _09731_ vssd1 vssd1 vccd1 vccd1 _09732_ sky130_fd_sc_hd__o21ai_2
XFILLER_70_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10636_ rbzero.tex_g1\[44\] rbzero.tex_g1\[45\] _03530_ vssd1 vssd1 vccd1 vccd1 _03538_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16143_ _07800_ _07712_ _08603_ vssd1 vssd1 vccd1 vccd1 _08755_ sky130_fd_sc_hd__or3_1
XFILLER_155_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13355_ _05793_ _05616_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__or2_1
XFILLER_122_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10567_ rbzero.tex_r0\[14\] rbzero.tex_r0\[13\] _03501_ vssd1 vssd1 vccd1 vccd1 _03502_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12306_ _04992_ rbzero.wall_tracer.trackDistX\[8\] rbzero.wall_tracer.trackDistX\[7\]
+ _04999_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__a22o_1
XFILLER_192_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16074_ _08527_ _08528_ vssd1 vssd1 vccd1 vccd1 _08687_ sky130_fd_sc_hd__nor2_1
XFILLER_155_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13286_ _05950_ _05974_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__xnor2_1
X_10498_ _03465_ vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__clkbuf_1
X_15025_ _07637_ _07638_ vssd1 vssd1 vccd1 vccd1 _07639_ sky130_fd_sc_hd__nand2_1
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19902_ _03112_ vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__clkinv_2
XFILLER_216_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12237_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__inv_2
XFILLER_68_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19833_ _03106_ vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__clkinv_2
XFILLER_190_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12168_ net33 vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__buf_2
XFILLER_111_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11119_ rbzero.traced_texVinit\[5\] rbzero.spi_registers.vshift\[2\] vssd1 vssd1
+ vccd1 vccd1 _03838_ sky130_fd_sc_hd__nand2_1
XFILLER_111_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19764_ _04632_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__inv_2
X_16976_ _09422_ _09383_ vssd1 vssd1 vccd1 vccd1 _09517_ sky130_fd_sc_hd__or2b_1
X_12099_ _04779_ _04805_ _04806_ _04793_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__a22o_1
XFILLER_232_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18715_ rbzero.wall_tracer.rayAddendY\[0\] _00013_ _02433_ _02441_ vssd1 vssd1 vccd1
+ vccd1 _00617_ sky130_fd_sc_hd__o22a_1
X_15927_ _07881_ _07885_ _08540_ vssd1 vssd1 vccd1 vccd1 _08541_ sky130_fd_sc_hd__a21o_1
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 i_gpout0_sel[3] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_6
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19695_ rbzero.pov.ready_buffer\[57\] _02963_ _03050_ vssd1 vssd1 vccd1 vccd1 _03051_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18646_ _02374_ _02377_ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__and2_1
X_15858_ _07814_ _07817_ vssd1 vssd1 vccd1 vccd1 _08472_ sky130_fd_sc_hd__nor2_1
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14809_ _07420_ _07421_ _07422_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__a21o_1
XFILLER_149_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18577_ _02308_ _02312_ _02317_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a21oi_1
XFILLER_224_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15789_ _08397_ _08401_ _08402_ vssd1 vssd1 vccd1 vccd1 _08403_ sky130_fd_sc_hd__a21oi_1
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17528_ _10062_ _10064_ vssd1 vssd1 vccd1 vccd1 _10065_ sky130_fd_sc_hd__or2_1
XFILLER_166_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17459_ _09994_ _09995_ _09996_ vssd1 vssd1 vccd1 vccd1 _09997_ sky130_fd_sc_hd__nand3_1
XFILLER_177_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20470_ net119 _00486_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19129_ rbzero.othery\[1\] _02723_ _02734_ _02728_ vssd1 vssd1 vccd1 vccd1 _00738_
+ sky130_fd_sc_hd__o211a_1
XFILLER_203_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21022_ net110 _01038_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20806_ _00024_ _00822_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20737_ net107 _00753_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11470_ rbzero.tex_r1\[1\] rbzero.tex_r1\[0\] _04168_ vssd1 vssd1 vccd1 vccd1 _04188_
+ sky130_fd_sc_hd__mux2_1
XFILLER_221_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20668_ net78 _00684_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10421_ _03423_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20599_ net82 _00615_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_104_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13140_ _05827_ _05828_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__xnor2_1
X_10352_ _03386_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13071_ _05650_ _05665_ _05759_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__a21bo_1
XFILLER_140_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10283_ _03350_ vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12022_ net8 net7 _04730_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__and3_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16830_ _09158_ _09121_ vssd1 vssd1 vccd1 vccd1 _09372_ sky130_fd_sc_hd__or2b_1
XFILLER_215_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13973_ _06609_ _06614_ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__xnor2_1
X_16761_ rbzero.wall_tracer.trackDistX\[-8\] rbzero.wall_tracer.stepDistX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _09311_ sky130_fd_sc_hd__nor2_1
XFILLER_120_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18500_ _02221_ _02233_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__nor2_1
X_15712_ _07470_ _07593_ _07971_ _08256_ vssd1 vssd1 vccd1 vccd1 _08326_ sky130_fd_sc_hd__o22ai_1
X_12924_ _05489_ _05612_ _05525_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__a21oi_4
XFILLER_111_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16692_ rbzero.traced_texa\[-4\] _09262_ _09263_ rbzero.wall_tracer.visualWallDist\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__a22o_1
X_19480_ _02907_ vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__clkbuf_1
XFILLER_234_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18431_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__nand2_1
X_15643_ _08256_ _07842_ vssd1 vssd1 vccd1 vccd1 _08257_ sky130_fd_sc_hd__nor2_1
X_12855_ _05481_ _05542_ _05543_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__o21ai_1
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11806_ rbzero.tex_b1\[49\] rbzero.tex_b1\[48\] _04032_ vssd1 vssd1 vccd1 vccd1 _04520_
+ sky130_fd_sc_hd__mux2_1
X_18362_ _02119_ _02120_ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__or2b_1
X_15574_ _08179_ _08185_ _08187_ vssd1 vssd1 vccd1 vccd1 _08188_ sky130_fd_sc_hd__a21oi_2
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12786_ _05438_ _05372_ _05375_ _05417_ _05462_ _05463_ vssd1 vssd1 vccd1 vccd1 _05475_
+ sky130_fd_sc_hd__mux4_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _08771_ _09607_ _09721_ _09722_ _09851_ vssd1 vssd1 vccd1 vccd1 _09852_ sky130_fd_sc_hd__a32oi_2
XFILLER_187_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14525_ _07177_ _07162_ _07201_ _07099_ vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__o211ai_4
XFILLER_159_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ rbzero.tex_b0\[58\] _03962_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__and2_1
X_18293_ _02058_ _02059_ _02060_ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__o21ai_1
XFILLER_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17244_ _09779_ _09781_ vssd1 vssd1 vccd1 vccd1 _09783_ sky130_fd_sc_hd__or2_1
X_14456_ _07141_ _07142_ _05527_ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__a21oi_1
XFILLER_147_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11668_ rbzero.tex_g1\[19\] rbzero.tex_g1\[18\] _04378_ vssd1 vssd1 vccd1 vccd1 _04384_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13407_ _06090_ _06091_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__or2_1
X_17175_ _09713_ _09714_ vssd1 vssd1 vccd1 vccd1 _09715_ sky130_fd_sc_hd__and2_1
XFILLER_200_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10619_ rbzero.tex_g1\[52\] rbzero.tex_g1\[53\] _03519_ vssd1 vssd1 vccd1 vccd1 _03529_
+ sky130_fd_sc_hd__mux2_1
X_14387_ _07028_ _07052_ _07063_ _07074_ _07075_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__a41o_1
XFILLER_155_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11599_ _03910_ _04313_ _04314_ _04315_ _03920_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__o221a_1
XFILLER_227_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16126_ _08730_ _08737_ vssd1 vssd1 vccd1 vccd1 _08738_ sky130_fd_sc_hd__xnor2_1
XFILLER_196_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13338_ _05995_ _06017_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16057_ _04937_ _07617_ vssd1 vssd1 vccd1 vccd1 _08670_ sky130_fd_sc_hd__or2_1
XFILLER_196_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13269_ _05616_ _05659_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__or2_1
XFILLER_142_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15008_ _07602_ _07621_ vssd1 vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__or2_1
XFILLER_130_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19816_ _03105_ vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__clkinv_2
XFILLER_233_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19747_ rbzero.pov.ready_buffer\[19\] _03069_ _03070_ _02191_ _02832_ vssd1 vssd1
+ vccd1 vccd1 _01020_ sky130_fd_sc_hd__o221a_1
X_16959_ _09118_ _09500_ vssd1 vssd1 vccd1 vccd1 _09501_ sky130_fd_sc_hd__xnor2_1
XFILLER_133_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19678_ rbzero.debug_overlay.playerY\[1\] _03032_ _03036_ vssd1 vssd1 vccd1 vccd1
+ _03037_ sky130_fd_sc_hd__a21o_1
XFILLER_237_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18629_ rbzero.debug_overlay.playerX\[3\] _02362_ _03797_ vssd1 vssd1 vccd1 vccd1
+ _02363_ sky130_fd_sc_hd__mux2_1
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_11 _07189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_22 rbzero.wall_tracer.visualWallDist\[-5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20522_ net113 _00538_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_33 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_44 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20453_ net117 _00004_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_193_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20384_ net131 _00415_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_84_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21005_ net56 _01021_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_247_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10970_ rbzero.tex_b0\[14\] rbzero.tex_b0\[13\] _03704_ vssd1 vssd1 vccd1 vccd1 _03713_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12640_ _05323_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__nor2_1
XFILLER_93_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12571_ _05258_ _05259_ _05219_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__mux2_2
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14310_ _06630_ _06998_ vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__and2_1
XFILLER_168_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11522_ _04226_ _04207_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__and2_2
X_15290_ _07873_ _07874_ _07903_ vssd1 vssd1 vccd1 vccd1 _07904_ sky130_fd_sc_hd__nand3_1
XFILLER_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14241_ _06921_ _06929_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__nand2_1
X_11453_ rbzero.tex_r1\[31\] _04142_ _04144_ _03929_ vssd1 vssd1 vccd1 vccd1 _04171_
+ sky130_fd_sc_hd__a31o_1
XFILLER_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10404_ _03414_ vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__clkbuf_1
X_14172_ _06859_ _06860_ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11384_ gpout0.vpos\[5\] _04102_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__or2_2
XFILLER_194_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13123_ _05809_ _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10335_ rbzero.tex_r1\[57\] rbzero.tex_r1\[58\] _03377_ vssd1 vssd1 vccd1 vccd1 _03378_
+ sky130_fd_sc_hd__mux2_1
X_18980_ rbzero.pov.spi_buffer\[38\] rbzero.pov.ready_buffer\[38\] _02640_ vssd1 vssd1
+ vccd1 vccd1 _02650_ sky130_fd_sc_hd__mux2_1
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17931_ _01498_ _01608_ _01607_ vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__a21oi_2
X_13054_ _05608_ _05619_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__nor2_1
XFILLER_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10266_ _03341_ vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12005_ net17 _04677_ _04701_ _04714_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__a31o_1
XFILLER_230_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17862_ _01627_ _01644_ vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__xnor2_2
XFILLER_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10197_ _03305_ vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19601_ _02727_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__buf_2
X_16813_ _09346_ _09348_ _09347_ vssd1 vssd1 vccd1 vccd1 _09357_ sky130_fd_sc_hd__a21boi_1
XFILLER_94_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17793_ _09968_ _09463_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__nor2_1
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19532_ rbzero.pov.spi_buffer\[61\] rbzero.pov.spi_buffer\[62\] _02932_ vssd1 vssd1
+ vccd1 vccd1 _02935_ sky130_fd_sc_hd__mux2_1
X_16744_ rbzero.wall_tracer.trackDistX\[-10\] rbzero.wall_tracer.stepDistX\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _09296_ sky130_fd_sc_hd__nor2_1
XFILLER_219_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13956_ _06435_ _06343_ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__nor2_1
XFILLER_235_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12907_ _05497_ _05554_ _05594_ _05595_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__o22a_1
X_19463_ _02898_ vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__clkbuf_1
X_13887_ _06553_ _06554_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__xor2_1
X_16675_ rbzero.row_render.size\[10\] _09260_ _07208_ _09261_ vssd1 vssd1 vccd1 vccd1
+ _00508_ sky130_fd_sc_hd__a22o_1
XFILLER_235_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18414_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__nand2_1
X_15626_ _07890_ vssd1 vssd1 vccd1 vccd1 _08240_ sky130_fd_sc_hd__buf_4
X_12838_ _05478_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__clkbuf_4
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19394_ _02862_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__buf_4
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18345_ _05002_ _02001_ _02106_ vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__a21oi_1
XFILLER_226_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12769_ _05360_ _05393_ _05397_ _05398_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__nand4_2
X_15557_ _08169_ _08170_ vssd1 vssd1 vccd1 vccd1 _08171_ sky130_fd_sc_hd__and2_2
XFILLER_148_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14508_ _07101_ _07187_ _07188_ vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__nand3_4
XFILLER_37_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18276_ rbzero.wall_tracer.trackDistY\[-4\] rbzero.wall_tracer.stepDistY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__nand2_1
X_15488_ _07992_ _08072_ vssd1 vssd1 vccd1 vccd1 _08102_ sky130_fd_sc_hd__and2_1
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17227_ rbzero.wall_tracer.trackDistX\[2\] rbzero.wall_tracer.stepDistX\[2\] vssd1
+ vssd1 vccd1 vccd1 _09767_ sky130_fd_sc_hd__or2_1
XFILLER_175_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput20 i_gpout2_sel[5] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_4
Xinput31 i_gpout4_sel[4] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_4
X_14439_ _07043_ _07034_ vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__nor2_1
XFILLER_239_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput42 i_reg_csb vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_8
XFILLER_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput53 i_vec_sclk vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_6
XFILLER_162_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17158_ _09575_ _09583_ _09582_ vssd1 vssd1 vccd1 vccd1 _09698_ sky130_fd_sc_hd__a21o_1
XFILLER_200_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16109_ _08719_ _08720_ vssd1 vssd1 vccd1 vccd1 _08721_ sky130_fd_sc_hd__nand2_1
XFILLER_143_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17089_ _09627_ _09629_ vssd1 vssd1 vccd1 vccd1 _09630_ sky130_fd_sc_hd__xor2_1
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20505_ net133 _00521_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20436_ net135 _00467_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20367_ _03287_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_7059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20298_ _03258_ vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__clkinv_2
XTAP_6347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13810_ _06457_ _06498_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__xnor2_1
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14790_ rbzero.debug_overlay.playerY\[-4\] rbzero.debug_overlay.playerY\[-5\] _07358_
+ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__or3_1
XFILLER_21_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13741_ _06418_ _06420_ _06429_ _06417_ _06405_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__o32ai_4
XFILLER_186_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10953_ _03604_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__clkbuf_4
XFILLER_21_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16460_ _09065_ _09066_ _09068_ vssd1 vssd1 vccd1 vccd1 _09070_ sky130_fd_sc_hd__a21o_1
XFILLER_231_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13672_ _06351_ _06360_ _06355_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__a21oi_1
XFILLER_243_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10884_ rbzero.tex_b0\[55\] rbzero.tex_b0\[54\] _03660_ vssd1 vssd1 vccd1 vccd1 _03668_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15411_ _08005_ _08022_ vssd1 vssd1 vccd1 vccd1 _08025_ sky130_fd_sc_hd__nor2_1
X_12623_ _05288_ _05311_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__nand2_1
X_16391_ _08997_ _09000_ vssd1 vssd1 vccd1 vccd1 _09001_ sky130_fd_sc_hd__xnor2_1
XFILLER_223_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18130_ _01908_ _01910_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__nor2_1
XFILLER_185_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15342_ _07588_ _07615_ _07639_ vssd1 vssd1 vccd1 vccd1 _07956_ sky130_fd_sc_hd__and3_1
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12554_ rbzero.wall_tracer.visualWallDist\[-7\] rbzero.wall_tracer.rcp_sel\[2\] vssd1
+ vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__or2_1
XFILLER_106_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11505_ _03780_ gpout0.hpos\[4\] _04215_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__nor3_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18061_ _01840_ _01841_ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__xnor2_1
X_15273_ _07878_ _07886_ _07884_ vssd1 vssd1 vccd1 vccd1 _07887_ sky130_fd_sc_hd__o21ai_1
XFILLER_185_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12485_ rbzero.debug_overlay.facingX\[-1\] rbzero.wall_tracer.rayAddendX\[7\] vssd1
+ vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__nand2_1
XFILLER_32_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17012_ _09547_ _09552_ vssd1 vssd1 vccd1 vccd1 _09553_ sky130_fd_sc_hd__and2_1
X_14224_ _06891_ _06912_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__nand2_1
XFILLER_156_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11436_ rbzero.tex_r1\[34\] _03925_ _03915_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__a21o_1
XFILLER_193_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14155_ _06137_ _06483_ vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__nor2_1
X_11367_ rbzero.row_render.size\[0\] gpout0.hpos\[1\] vssd1 vssd1 vccd1 vccd1 _04086_
+ sky130_fd_sc_hd__or2_1
XFILLER_193_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13106_ _05608_ _05660_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__or2_1
XFILLER_98_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10318_ rbzero.tex_b1\[1\] rbzero.tex_b1\[2\] _03366_ vssd1 vssd1 vccd1 vccd1 _03369_
+ sky130_fd_sc_hd__mux2_1
X_14086_ _06757_ _06773_ _06774_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__a21bo_1
XFILLER_119_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18963_ _02641_ vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__clkbuf_1
X_11298_ _04007_ _04010_ _04016_ _03950_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__a211o_1
XFILLER_234_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17914_ _01695_ _01696_ vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__or2_1
X_13037_ _05706_ _05707_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__and2_1
X_10249_ _03332_ vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18894_ _02602_ _02589_ _02603_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__and3b_1
XFILLER_67_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17845_ _10111_ _01587_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__nand2_1
XFILLER_227_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17776_ _01556_ _01558_ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__nand2_1
XFILLER_81_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14988_ _07599_ _07601_ vssd1 vssd1 vccd1 vccd1 _07602_ sky130_fd_sc_hd__and2_2
XFILLER_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19515_ rbzero.pov.spi_buffer\[53\] rbzero.pov.spi_buffer\[54\] _02921_ vssd1 vssd1
+ vccd1 vccd1 _02926_ sky130_fd_sc_hd__mux2_1
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16727_ rbzero.wall_tracer.trackDistX\[-12\] rbzero.wall_tracer.stepDistX\[-12\]
+ vssd1 vssd1 vccd1 vccd1 _09281_ sky130_fd_sc_hd__or2_1
X_13939_ _06575_ _06627_ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__nor2_1
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19446_ rbzero.pov.spi_buffer\[20\] rbzero.pov.spi_buffer\[21\] _02888_ vssd1 vssd1
+ vccd1 vccd1 _02890_ sky130_fd_sc_hd__mux2_1
X_16658_ _03728_ vssd1 vssd1 vccd1 vccd1 _09256_ sky130_fd_sc_hd__buf_4
XFILLER_126_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15609_ _08222_ vssd1 vssd1 vccd1 vccd1 _08223_ sky130_fd_sc_hd__clkbuf_4
X_19377_ _02860_ vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__clkinv_2
XFILLER_72_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16589_ _07243_ vssd1 vssd1 vccd1 vccd1 _09198_ sky130_fd_sc_hd__inv_2
XFILLER_245_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18328_ _02089_ _02090_ _02091_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__a21o_1
XFILLER_176_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18259_ rbzero.wall_tracer.trackDistY\[-7\] _01996_ _02032_ _09317_ vssd1 vssd1 vccd1
+ vccd1 _00570_ sky130_fd_sc_hd__o22a_1
XFILLER_50_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21270_ _00319_ _01286_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20221_ _03236_ _03238_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20152_ _03177_ _03178_ _03179_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__nand3_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20083_ _03131_ vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__clkinv_2
XFILLER_44_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20985_ net65 _01001_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _04962_ rbzero.wall_tracer.trackDistY\[-7\] rbzero.wall_tracer.trackDistY\[-8\]
+ _04963_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__a22o_1
XFILLER_138_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11221_ _03901_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__clkbuf_4
XFILLER_107_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20419_ net128 _00450_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21399_ net83 _01415_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11152_ _03870_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__inv_2
XTAP_6111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15960_ rbzero.debug_overlay.playerY\[-8\] vssd1 vssd1 vccd1 vccd1 _08574_ sky130_fd_sc_hd__inv_2
X_11083_ _03805_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14911_ rbzero.wall_tracer.stepDistY\[-11\] vssd1 vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__inv_2
XFILLER_118_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15891_ _07859_ _07867_ _08504_ vssd1 vssd1 vccd1 vccd1 _08505_ sky130_fd_sc_hd__a21bo_1
XTAP_5465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17630_ _09684_ _09022_ _08850_ _08978_ vssd1 vssd1 vccd1 vccd1 _10166_ sky130_fd_sc_hd__or4_1
XTAP_5498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ _07435_ _07442_ _07443_ _07455_ vssd1 vssd1 vccd1 vccd1 _07456_ sky130_fd_sc_hd__or4_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17561_ _07631_ _09955_ vssd1 vssd1 vccd1 vccd1 _10098_ sky130_fd_sc_hd__nor2_1
X_14773_ _07384_ _07385_ _07386_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__a21o_2
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11985_ net19 net20 vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__and2b_1
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19300_ rbzero.pov.spi_done rbzero.pov.ready _02832_ _02836_ vssd1 vssd1 vccd1 vccd1
+ _00807_ sky130_fd_sc_hd__o211a_1
XFILLER_229_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16512_ _08994_ _09008_ _09006_ vssd1 vssd1 vccd1 vccd1 _09121_ sky130_fd_sc_hd__a21o_1
XFILLER_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13724_ _06326_ _06411_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__xor2_1
XFILLER_182_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10936_ _03695_ vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17492_ _07291_ _09283_ _10029_ vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19231_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.new_floor\[2\]
+ _02795_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__mux2_1
XFILLER_108_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16443_ _09048_ _09052_ vssd1 vssd1 vccd1 vccd1 _09053_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13655_ _05861_ _06343_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__nor2_1
X_10867_ rbzero.tex_b0\[63\] rbzero.tex_b0\[62\] _03649_ vssd1 vssd1 vccd1 vccd1 _03659_
+ sky130_fd_sc_hd__mux2_1
XFILLER_220_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12606_ _05220_ _05294_ _05280_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__a21o_1
XFILLER_9_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19162_ _02742_ _02755_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__and2_1
X_16374_ _07519_ _08663_ vssd1 vssd1 vccd1 vccd1 _08984_ sky130_fd_sc_hd__or2_1
X_13586_ _06273_ _06274_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__nand2_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ rbzero.tex_g0\[32\] rbzero.tex_g0\[31\] _03616_ vssd1 vssd1 vccd1 vccd1 _03623_
+ sky130_fd_sc_hd__mux2_1
XFILLER_223_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18113_ _01760_ _01795_ _01893_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a21bo_1
XFILLER_157_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15325_ _07664_ _07709_ vssd1 vssd1 vccd1 vccd1 _07939_ sky130_fd_sc_hd__nor2_1
X_12537_ _05167_ _05225_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__xnor2_2
XFILLER_9_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19093_ _02710_ vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18044_ _01722_ _01725_ _01723_ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__o21ai_1
XFILLER_157_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15256_ _07856_ _07857_ _07868_ vssd1 vssd1 vccd1 vccd1 _07870_ sky130_fd_sc_hd__a21o_1
XFILLER_173_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12468_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__or2_1
XFILLER_173_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14207_ _06895_ _06892_ vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__xnor2_1
X_11419_ rbzero.tex_r1\[46\] _04013_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__and2_1
X_15187_ _07388_ _07552_ _07800_ _07424_ vssd1 vssd1 vccd1 vccd1 _07801_ sky130_fd_sc_hd__o22ai_1
X_12399_ _05042_ _05038_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__or2b_1
XFILLER_235_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14138_ _06742_ _06826_ vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__nand2_1
XFILLER_158_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19995_ _03122_ vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__clkinv_2
XFILLER_154_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14069_ _06724_ _06716_ _06723_ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__nand3_1
X_18946_ _02632_ vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18877_ rbzero.spi_registers.spi_counter\[1\] rbzero.spi_registers.spi_counter\[0\]
+ _02576_ vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__nand3_1
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17828_ _03797_ _01610_ _01611_ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__or3_1
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17759_ _01539_ _01541_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__nand2_1
XFILLER_70_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20770_ net103 _00786_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19429_ rbzero.pov.spi_buffer\[12\] rbzero.pov.spi_buffer\[13\] _02877_ vssd1 vssd1
+ vccd1 vccd1 _02881_ sky130_fd_sc_hd__mux2_1
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21322_ _00345_ _01338_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21253_ _00302_ _01269_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20204_ _03223_ _03224_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__xnor2_1
XFILLER_116_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21184_ _00233_ _01200_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20135_ _03163_ _03164_ _03165_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__o21ai_1
XFILLER_213_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20066_ _03129_ vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__clkinv_2
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11770_ rbzero.tex_b0\[29\] rbzero.tex_b0\[28\] _04001_ vssd1 vssd1 vccd1 vccd1 _04485_
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20968_ net71 _00984_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _03582_ vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20899_ net60 _00915_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13440_ _05488_ _05625_ vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__nand2_1
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10652_ _03546_ vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13371_ _06027_ _06059_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__or2_1
XFILLER_210_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10583_ rbzero.tex_r0\[6\] rbzero.tex_r0\[5\] _03501_ vssd1 vssd1 vccd1 vccd1 _03510_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15110_ _07716_ _07723_ vssd1 vssd1 vccd1 vccd1 _07724_ sky130_fd_sc_hd__xor2_1
X_12322_ rbzero.wall_tracer.trackDistY\[-8\] vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__inv_2
X_16090_ _08700_ _08701_ vssd1 vssd1 vccd1 vccd1 _08703_ sky130_fd_sc_hd__and2_1
XFILLER_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15041_ _07100_ _07210_ vssd1 vssd1 vccd1 vccd1 _07655_ sky130_fd_sc_hd__and2_1
XFILLER_68_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12253_ rbzero.wall_tracer.trackDistX\[-3\] vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__inv_2
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11204_ _03920_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__buf_4
XFILLER_68_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12184_ _04883_ o_rgb[14] vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__or2_1
XFILLER_122_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18800_ _02509_ _04260_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__nand2_1
XFILLER_150_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11135_ _03850_ _03849_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__nand2_1
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19780_ _04631_ _03085_ _03086_ _03031_ vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__o211a_1
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16992_ _09531_ _09532_ vssd1 vssd1 vccd1 vccd1 _09533_ sky130_fd_sc_hd__nand2_1
XFILLER_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18731_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__or2_1
X_15943_ _08555_ _08556_ vssd1 vssd1 vccd1 vccd1 _08557_ sky130_fd_sc_hd__xnor2_1
XTAP_5240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11066_ rbzero.wall_tracer.state\[8\] vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__inv_2
XFILLER_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18662_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__or2_1
XFILLER_92_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15874_ _07824_ _07847_ _08486_ _08487_ vssd1 vssd1 vccd1 vccd1 _08488_ sky130_fd_sc_hd__or4bb_1
XTAP_5295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17613_ _07294_ _09283_ _10149_ vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__a21oi_1
XFILLER_149_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14825_ _07436_ _07438_ rbzero.wall_tracer.state\[13\] vssd1 vssd1 vccd1 vccd1 _07439_
+ sky130_fd_sc_hd__a21o_1
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18593_ rbzero.debug_overlay.vplaneX\[0\] _02191_ _02318_ _02275_ vssd1 vssd1 vccd1
+ vccd1 _02333_ sky130_fd_sc_hd__a211oi_1
XFILLER_221_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ _09939_ _09934_ vssd1 vssd1 vccd1 vccd1 _10081_ sky130_fd_sc_hd__and2b_1
XFILLER_233_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14756_ _05236_ _05247_ _05242_ _07369_ vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__or4_1
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11968_ _03288_ _04592_ _04631_ _04632_ net15 _04671_ vssd1 vssd1 vccd1 vccd1 _04678_
+ sky130_fd_sc_hd__mux4_1
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13707_ _06353_ _06354_ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17475_ _09788_ _09877_ _10012_ vssd1 vssd1 vccd1 vccd1 _10013_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10919_ _03686_ vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14687_ rbzero.wall_tracer.stepDistX\[-2\] _07196_ _07316_ vssd1 vssd1 vccd1 vccd1
+ _07318_ sky130_fd_sc_hd__mux2_1
X_11899_ net73 vssd1 vssd1 vccd1 vccd1 o_tex_sclk sky130_fd_sc_hd__inv_2
XFILLER_220_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19214_ _02788_ vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16426_ _08915_ _08925_ _08924_ vssd1 vssd1 vccd1 vccd1 _09036_ sky130_fd_sc_hd__o21bai_1
XFILLER_34_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13638_ _06314_ _06326_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__xor2_2
XFILLER_220_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19145_ rbzero.spi_registers.new_leak\[0\] _02745_ vssd1 vssd1 vccd1 vccd1 _02746_
+ sky130_fd_sc_hd__or2_1
XFILLER_201_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16357_ _08961_ _08959_ vssd1 vssd1 vccd1 vccd1 _08967_ sky130_fd_sc_hd__and2b_1
X_13569_ _06256_ _06257_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__nor2_1
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15308_ _07623_ _07628_ vssd1 vssd1 vccd1 vccd1 _07922_ sky130_fd_sc_hd__and2b_1
XFILLER_145_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19076_ _02700_ vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__clkbuf_1
X_16288_ _07742_ _08760_ _08757_ _08755_ vssd1 vssd1 vccd1 vccd1 _08899_ sky130_fd_sc_hd__o31a_1
XFILLER_172_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18027_ _01802_ _01803_ _01807_ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__and3_1
XFILLER_161_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15239_ _07850_ _07851_ _07830_ vssd1 vssd1 vccd1 vccd1 _07853_ sky130_fd_sc_hd__a21o_1
XFILLER_161_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19978_ _03120_ vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__clkinv_2
XFILLER_99_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18929_ _02623_ vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20822_ _00040_ _00838_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20753_ net105 _00769_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20684_ net75 _00700_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[64\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21305_ net129 _01321_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_237_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21236_ _00285_ _01252_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21167_ _00216_ _01183_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20118_ rbzero.texV\[-9\] _02989_ _03142_ _03152_ vssd1 vssd1 vccd1 vccd1 _01309_
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21098_ _00147_ _01114_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12940_ _05628_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__buf_2
XFILLER_4_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20049_ _03128_ vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__clkinv_2
XFILLER_86_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _05506_ _05418_ _05430_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__mux2_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ rbzero.wall_tracer.trackDistX\[-6\] rbzero.wall_tracer.trackDistY\[-6\] _07258_
+ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__mux2_1
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11822_ rbzero.tex_b1\[45\] rbzero.tex_b1\[44\] _03903_ vssd1 vssd1 vccd1 vccd1 _04536_
+ sky130_fd_sc_hd__mux2_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _08199_ _08200_ vssd1 vssd1 vccd1 vccd1 _08204_ sky130_fd_sc_hd__nor2_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14541_ _05440_ _07007_ vssd1 vssd1 vccd1 vccd1 _07214_ sky130_fd_sc_hd__nand2_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11753_ rbzero.tex_b0\[43\] rbzero.tex_b0\[42\] _04001_ vssd1 vssd1 vccd1 vccd1 _04468_
+ sky130_fd_sc_hd__mux2_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10704_ _03573_ vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__clkbuf_1
X_17260_ _09684_ _09022_ _08718_ _08985_ vssd1 vssd1 vccd1 vccd1 _09799_ sky130_fd_sc_hd__or4_1
XFILLER_144_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14472_ rbzero.wall_tracer.stepDistY\[-9\] _07157_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _07158_ sky130_fd_sc_hd__mux2_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ rbzero.tex_g1\[15\] rbzero.tex_g1\[14\] _03980_ vssd1 vssd1 vccd1 vccd1 _04400_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16211_ _08691_ _08692_ _08689_ vssd1 vssd1 vccd1 vccd1 _08823_ sky130_fd_sc_hd__o21a_1
X_13423_ _06106_ _06110_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__nor2_1
X_10635_ _03537_ vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__clkbuf_1
X_17191_ _04938_ rbzero.wall_tracer.stepDistX\[11\] vssd1 vssd1 vccd1 vccd1 _09731_
+ sky130_fd_sc_hd__nand2_2
XFILLER_186_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16142_ _08752_ _08753_ vssd1 vssd1 vccd1 vccd1 _08754_ sky130_fd_sc_hd__xnor2_1
X_13354_ _05635_ _05660_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__or2_1
XFILLER_154_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10566_ _03445_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__clkbuf_4
X_12305_ rbzero.wall_tracer.trackDistY\[7\] vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__inv_2
XFILLER_182_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16073_ _08658_ _08685_ vssd1 vssd1 vccd1 vccd1 _08686_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13285_ _05951_ _05972_ _05973_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__a21oi_1
X_10497_ rbzero.tex_r0\[47\] rbzero.tex_r0\[46\] _03457_ vssd1 vssd1 vccd1 vccd1 _03465_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15024_ _07630_ _07636_ vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__or2_1
XFILLER_170_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12236_ _04931_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__buf_4
X_19901_ _03112_ vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__clkinv_2
XFILLER_155_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19832_ _03106_ vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__clkinv_2
X_12167_ net34 vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__buf_2
XFILLER_155_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11118_ rbzero.traced_texVinit\[5\] rbzero.spi_registers.vshift\[2\] vssd1 vssd1
+ vccd1 vccd1 _03837_ sky130_fd_sc_hd__or2_1
X_19763_ _03072_ vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__clkbuf_1
X_16975_ _09371_ _09381_ _09379_ vssd1 vssd1 vccd1 vccd1 _09516_ sky130_fd_sc_hd__a21o_1
XFILLER_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12098_ net49 net40 net39 net41 _04773_ _04768_ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__mux4_1
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18714_ _02166_ _02439_ _02440_ _09254_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__a31o_1
XFILLER_232_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15926_ _08538_ _08539_ vssd1 vssd1 vccd1 vccd1 _08540_ sky130_fd_sc_hd__xor2_1
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ _03765_ _03768_ _03775_ _03776_ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__and4b_1
XFILLER_237_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19694_ _02833_ _03049_ _03012_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__o21a_1
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput7 i_gpout0_sel[4] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_4
XFILLER_225_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18645_ _02375_ _02376_ _02374_ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__nand3b_1
XFILLER_225_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15857_ _08461_ _08470_ vssd1 vssd1 vccd1 vccd1 _08471_ sky130_fd_sc_hd__xor2_1
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14808_ _04927_ rbzero.wall_tracer.stepDistX\[-6\] vssd1 vssd1 vccd1 vccd1 _07422_
+ sky130_fd_sc_hd__nor2_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18576_ rbzero.debug_overlay.vplaneX\[0\] _02305_ _02316_ vssd1 vssd1 vccd1 vccd1
+ _02317_ sky130_fd_sc_hd__a21o_1
X_15788_ _08392_ _08396_ vssd1 vssd1 vccd1 vccd1 _08402_ sky130_fd_sc_hd__nor2_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17527_ _09022_ _08724_ _09922_ _10063_ vssd1 vssd1 vccd1 vccd1 _10064_ sky130_fd_sc_hd__o31a_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14739_ _07351_ rbzero.wall_tracer.stepDistY\[-4\] _07352_ vssd1 vssd1 vccd1 vccd1
+ _07353_ sky130_fd_sc_hd__a21oi_2
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17458_ _09856_ _09864_ _09863_ vssd1 vssd1 vccd1 vccd1 _09996_ sky130_fd_sc_hd__a21o_1
XFILLER_221_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16409_ _07591_ _07736_ _07520_ _09018_ vssd1 vssd1 vccd1 vccd1 _09019_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_203_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17389_ _09925_ _09926_ vssd1 vssd1 vccd1 vccd1 _09927_ sky130_fd_sc_hd__or2_1
XFILLER_20_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19128_ rbzero.spi_registers.new_other\[1\] _02725_ vssd1 vssd1 vccd1 vccd1 _02734_
+ sky130_fd_sc_hd__or2_1
XFILLER_185_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19059_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.spi_buffer\[0\]
+ _02690_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__mux2_1
XFILLER_133_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21021_ net110 _01037_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20805_ _00023_ _00821_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20736_ net105 _00752_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20667_ net68 _00683_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10420_ rbzero.tex_r1\[17\] rbzero.tex_r1\[18\] _03422_ vssd1 vssd1 vccd1 vccd1 _03423_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20598_ net82 _00614_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_109_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10351_ rbzero.tex_r1\[49\] rbzero.tex_r1\[50\] _03377_ vssd1 vssd1 vccd1 vccd1 _03386_
+ sky130_fd_sc_hd__mux2_1
XFILLER_104_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13070_ _05656_ _05664_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__or2b_1
X_10282_ rbzero.tex_b1\[18\] rbzero.tex_b1\[19\] _03344_ vssd1 vssd1 vccd1 vccd1 _03350_
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12021_ net4 net5 net6 vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__a21o_1
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21219_ _00268_ _01235_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16760_ _09279_ _08573_ vssd1 vssd1 vccd1 vccd1 _09310_ sky130_fd_sc_hd__nor2_1
XFILLER_76_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13972_ _06655_ _06660_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__nor2_1
XFILLER_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15711_ _07467_ _07986_ vssd1 vssd1 vccd1 vccd1 _08325_ sky130_fd_sc_hd__or2_1
XFILLER_247_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12923_ _05512_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__clkbuf_4
XFILLER_20_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16691_ rbzero.traced_texa\[-5\] _09262_ _09263_ rbzero.wall_tracer.visualWallDist\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__a22o_1
XFILLER_111_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18430_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__or2_1
X_15642_ _07420_ _07421_ vssd1 vssd1 vccd1 vccd1 _08256_ sky130_fd_sc_hd__and2_2
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _05527_ _05486_ _05467_ _05538_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__a22o_1
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18361_ rbzero.wall_tracer.trackDistY\[8\] rbzero.wall_tracer.stepDistY\[8\] vssd1
+ vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__nand2_1
XFILLER_203_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11805_ _04519_ vssd1 vssd1 vccd1 vccd1 o_rgb[22] sky130_fd_sc_hd__inv_2
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15573_ _08157_ _08186_ vssd1 vssd1 vccd1 vccd1 _08187_ sky130_fd_sc_hd__or2_1
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _05360_ _05473_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__or2_2
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _08923_ _09470_ _08272_ vssd1 vssd1 vccd1 vccd1 _09851_ sky130_fd_sc_hd__a21o_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14524_ _07133_ _07063_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__or2_1
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18292_ _02058_ _02059_ _02060_ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__or3_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11736_ rbzero.tex_b0\[57\] rbzero.tex_b0\[56\] _04013_ vssd1 vssd1 vccd1 vccd1 _04451_
+ sky130_fd_sc_hd__mux2_1
XFILLER_202_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17243_ _09779_ _09781_ vssd1 vssd1 vccd1 vccd1 _09782_ sky130_fd_sc_hd__nand2_1
XFILLER_41_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14455_ _07105_ _07103_ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__nand2_1
XFILLER_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11667_ _03994_ _04377_ _04382_ _03956_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__a211o_1
X_13406_ _06094_ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__inv_2
X_17174_ _09705_ _09712_ vssd1 vssd1 vccd1 vccd1 _09714_ sky130_fd_sc_hd__or2_1
XFILLER_122_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10618_ _03528_ vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__clkbuf_1
X_14386_ _05440_ _05405_ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__or2_2
XFILLER_167_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11598_ rbzero.tex_g0\[31\] _03938_ _03940_ _03915_ vssd1 vssd1 vccd1 vccd1 _04315_
+ sky130_fd_sc_hd__a31o_1
X_16125_ _08734_ _08736_ vssd1 vssd1 vccd1 vccd1 _08737_ sky130_fd_sc_hd__xor2_1
XFILLER_183_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13337_ _05981_ _06022_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__xor2_1
XFILLER_143_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10549_ _03492_ vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16056_ _07792_ _08668_ vssd1 vssd1 vccd1 vccd1 _08669_ sky130_fd_sc_hd__or2_1
XFILLER_170_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13268_ _05564_ _05672_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__or2_1
XFILLER_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15007_ _07620_ vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__buf_2
X_12219_ o_vsync rbzero.wall_tracer.state\[2\] _04920_ vssd1 vssd1 vccd1 vccd1 _04922_
+ sky130_fd_sc_hd__and3_1
XFILLER_97_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13199_ _05564_ _05622_ _05886_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__or3b_1
XFILLER_243_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19815_ _02862_ vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__buf_4
XFILLER_96_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16958_ _09497_ _09499_ vssd1 vssd1 vccd1 vccd1 _09500_ sky130_fd_sc_hd__xor2_1
XFILLER_110_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19746_ rbzero.pov.ready_buffer\[18\] _03067_ _03068_ rbzero.debug_overlay.vplaneX\[-2\]
+ _03015_ vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__a221o_1
XFILLER_244_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15909_ _08505_ _08522_ vssd1 vssd1 vccd1 vccd1 _08523_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19677_ rbzero.debug_overlay.playerY\[1\] _03032_ _02962_ vssd1 vssd1 vccd1 vccd1
+ _03036_ sky130_fd_sc_hd__o21ai_1
X_16889_ _09427_ _09430_ vssd1 vssd1 vccd1 vccd1 _09431_ sky130_fd_sc_hd__nand2_1
XFILLER_38_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18628_ _02360_ _02361_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18559_ _02279_ _02273_ _02288_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__nor3_1
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_12 _07840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_23 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20521_ net113 _00537_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_34 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_45 net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20452_ net118 _00003_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20383_ net121 _00414_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21004_ net82 _01020_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12570_ rbzero.wall_tracer.visualWallDist\[-9\] _05096_ rbzero.wall_tracer.rcp_sel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__mux2_1
XFILLER_19_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11521_ rbzero.debug_overlay.facingX\[-6\] _04237_ _04238_ rbzero.debug_overlay.facingX\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__a22o_1
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20719_ net88 _00735_ vssd1 vssd1 vccd1 vccd1 rbzero.otherx\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14240_ _06927_ _06928_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__and2_1
X_11452_ rbzero.tex_r1\[30\] _03961_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__and2_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10403_ rbzero.tex_r1\[25\] rbzero.tex_r1\[26\] _03411_ vssd1 vssd1 vccd1 vccd1 _03414_
+ sky130_fd_sc_hd__mux2_1
X_14171_ _06101_ _06482_ vssd1 vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__nor2_1
X_11383_ gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__inv_2
XFILLER_165_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13122_ _05693_ _05810_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__and2_1
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10334_ _03299_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__clkbuf_4
XFILLER_194_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17930_ _01711_ _01712_ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__and2_1
X_13053_ _05739_ _05741_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__or2_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ rbzero.tex_b1\[26\] rbzero.tex_b1\[27\] _03333_ vssd1 vssd1 vccd1 vccd1 _03341_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12004_ _04668_ _04705_ _04695_ _04713_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_78_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17861_ _01629_ _01643_ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10196_ rbzero.tex_b1\[59\] rbzero.tex_b1\[60\] _03300_ vssd1 vssd1 vccd1 vccd1 _03305_
+ sky130_fd_sc_hd__mux2_1
XFILLER_239_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16812_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.stepDistX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _09356_ sky130_fd_sc_hd__and2_1
X_19600_ _07493_ _02960_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__nand2_1
XFILLER_78_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17792_ _01458_ _01574_ _01575_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__o21ai_1
XFILLER_226_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19531_ _02934_ vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16743_ _09288_ _09289_ vssd1 vssd1 vccd1 vccd1 _09295_ sky130_fd_sc_hd__and2_1
XFILLER_207_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13955_ _06028_ _06305_ _06643_ vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__a21o_1
XFILLER_47_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12906_ _05412_ _05431_ _05497_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__o21ai_1
X_19462_ rbzero.pov.spi_buffer\[28\] rbzero.pov.spi_buffer\[29\] _02888_ vssd1 vssd1
+ vccd1 vccd1 _02898_ sky130_fd_sc_hd__mux2_1
XFILLER_228_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16674_ _09257_ vssd1 vssd1 vccd1 vccd1 _09261_ sky130_fd_sc_hd__buf_4
XFILLER_59_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13886_ _06559_ _06557_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__xor2_1
X_18413_ _09256_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__clkbuf_4
X_15625_ _08237_ _08238_ vssd1 vssd1 vccd1 vccd1 _08239_ sky130_fd_sc_hd__and2_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _05489_ _05512_ _05525_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__a21o_2
XFILLER_37_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19393_ _04702_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__buf_4
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _09351_ _02104_ _02105_ _10148_ _01995_ vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__o311a_1
XFILLER_199_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15556_ _08111_ _08168_ vssd1 vssd1 vccd1 vccd1 _08170_ sky130_fd_sc_hd__or2_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12768_ _05455_ _05456_ _05453_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__mux2_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _07133_ _07089_ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__or2_1
XFILLER_175_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18275_ rbzero.wall_tracer.trackDistY\[-4\] rbzero.wall_tracer.stepDistY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__nor2_1
XFILLER_147_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11719_ rbzero.tex_g1\[37\] rbzero.tex_g1\[36\] _03980_ vssd1 vssd1 vccd1 vccd1 _04435_
+ sky130_fd_sc_hd__mux2_1
X_15487_ _08075_ _08100_ vssd1 vssd1 vccd1 vccd1 _08101_ sky130_fd_sc_hd__nand2_1
XFILLER_148_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12699_ _05351_ _05354_ _05386_ _05387_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__or4_1
XFILLER_238_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17226_ rbzero.wall_tracer.trackDistX\[2\] rbzero.wall_tracer.stepDistX\[2\] vssd1
+ vssd1 vccd1 vccd1 _09766_ sky130_fd_sc_hd__nand2_1
XFILLER_200_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14438_ _07105_ _07125_ vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__or2_1
XFILLER_147_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput10 i_gpout1_sel[1] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_4
Xinput21 i_gpout3_sel[0] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_4
XFILLER_163_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput32 i_gpout4_sel[5] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_4
XFILLER_200_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput43 i_reg_mosi vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_6
XFILLER_239_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17157_ _09661_ _09696_ vssd1 vssd1 vccd1 vccd1 _09697_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14369_ _05593_ _07024_ vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__or2_1
XFILLER_171_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16108_ _07788_ _08718_ _08663_ _08429_ vssd1 vssd1 vccd1 vccd1 _08720_ sky130_fd_sc_hd__o22ai_1
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17088_ _09423_ _09492_ _09628_ vssd1 vssd1 vccd1 vccd1 _09629_ sky130_fd_sc_hd__a21boi_1
XFILLER_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16039_ _08650_ _08651_ vssd1 vssd1 vccd1 vccd1 _08652_ sky130_fd_sc_hd__xor2_1
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19729_ rbzero.pov.ready_buffer\[27\] _03061_ _03063_ rbzero.debug_overlay.facingY\[-4\]
+ _03066_ vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__a221o_1
XFILLER_244_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20504_ net132 _00520_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20435_ net135 _00466_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20366_ _02727_ _03285_ _03286_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__and3_1
XTAP_7016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20297_ _03258_ vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__clkinv_2
XTAP_6326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13740_ _06424_ _06427_ _06428_ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__o21a_1
XFILLER_112_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10952_ _03703_ vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13671_ _06355_ _06359_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__nor2_1
XFILLER_147_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10883_ _03667_ vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15410_ _07998_ _07982_ vssd1 vssd1 vccd1 vccd1 _08024_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12622_ _05220_ _05283_ _05280_ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__a21oi_2
XPHY_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16390_ _08998_ _08999_ vssd1 vssd1 vccd1 vccd1 _09000_ sky130_fd_sc_hd__and2b_1
XPHY_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15341_ _07931_ _07954_ vssd1 vssd1 vccd1 vccd1 _07955_ sky130_fd_sc_hd__xor2_1
XFILLER_129_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12553_ _05240_ _05241_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__xnor2_4
XPHY_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18060_ _07631_ _08787_ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__nor2_1
XFILLER_157_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11504_ _03803_ _04200_ _04217_ _04221_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__a211o_1
X_15272_ _07598_ vssd1 vssd1 vccd1 vccd1 _07886_ sky130_fd_sc_hd__clkbuf_4
XFILLER_145_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12484_ _05172_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__inv_2
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17011_ _09550_ _09551_ vssd1 vssd1 vccd1 vccd1 _09552_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14223_ _05668_ _06175_ _06421_ _06890_ vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__a31o_1
XFILLER_123_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11435_ rbzero.tex_r1\[35\] _03938_ _03940_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__and3_1
XFILLER_208_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14154_ _06811_ _06842_ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__xor2_1
XFILLER_197_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11366_ gpout0.hpos\[1\] gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__and2_1
XFILLER_99_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13105_ _05793_ _05621_ _05658_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__nor3_1
XFILLER_158_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10317_ _03368_ vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14085_ _06758_ _06759_ _06772_ vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__nand3_1
X_18962_ rbzero.pov.spi_buffer\[29\] rbzero.pov.ready_buffer\[29\] _02640_ vssd1 vssd1
+ vccd1 vccd1 _02641_ sky130_fd_sc_hd__mux2_1
X_11297_ _03932_ _04011_ _04012_ _04015_ _03946_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__o221a_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17913_ _01542_ _01545_ _01694_ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__and3_1
X_13036_ _05525_ _05700_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__nand2_1
X_10248_ rbzero.tex_b1\[34\] rbzero.tex_b1\[35\] _03322_ vssd1 vssd1 vccd1 vccd1 _03332_
+ sky130_fd_sc_hd__mux2_1
X_18893_ rbzero.spi_registers.spi_counter\[4\] rbzero.spi_registers.spi_counter\[3\]
+ _02594_ rbzero.spi_registers.spi_counter\[5\] vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a31o_1
XTAP_6860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17844_ _01573_ _01580_ _01626_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__a21o_1
XFILLER_113_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10179_ net46 net45 vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__xor2_4
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17775_ _01556_ _01558_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__nor2_1
XFILLER_130_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14987_ _07346_ _07600_ _07349_ vssd1 vssd1 vccd1 vccd1 _07601_ sky130_fd_sc_hd__a21oi_2
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16726_ rbzero.wall_tracer.trackDistX\[-12\] rbzero.wall_tracer.stepDistX\[-12\]
+ vssd1 vssd1 vccd1 vccd1 _09280_ sky130_fd_sc_hd__nand2_1
X_19514_ _02925_ vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__clkbuf_1
X_13938_ _06576_ _06622_ _06626_ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__o21a_1
XFILLER_130_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19445_ _02889_ vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__clkbuf_1
XFILLER_228_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16657_ _09254_ vssd1 vssd1 vccd1 vccd1 _09255_ sky130_fd_sc_hd__buf_2
X_13869_ _05434_ _06550_ _06548_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__o21ai_1
XFILLER_90_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15608_ _07350_ _07353_ vssd1 vssd1 vccd1 vccd1 _08222_ sky130_fd_sc_hd__and2_1
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19376_ _02860_ vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__clkinv_2
XFILLER_76_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16588_ _04939_ rbzero.wall_tracer.stepDistX\[7\] _08634_ vssd1 vssd1 vccd1 vccd1
+ _09197_ sky130_fd_sc_hd__a21boi_4
XFILLER_241_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18327_ _02082_ _02086_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__nand2_1
X_15539_ _07566_ _08060_ vssd1 vssd1 vccd1 vccd1 _08153_ sky130_fd_sc_hd__nor2_1
XFILLER_163_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18258_ _01997_ _02030_ _02031_ _02013_ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__a31o_1
XFILLER_191_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17209_ _09623_ _09625_ vssd1 vssd1 vccd1 vccd1 _09749_ sky130_fd_sc_hd__nor2_1
XFILLER_129_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18189_ _08918_ _08921_ _07886_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a21oi_2
XFILLER_129_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20220_ rbzero.traced_texa\[7\] rbzero.texV\[7\] _03237_ vssd1 vssd1 vccd1 vccd1
+ _03238_ sky130_fd_sc_hd__o21ai_1
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20151_ _03177_ _03178_ _03179_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__a21o_1
XFILLER_103_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20082_ _03131_ vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__clkinv_2
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20984_ net65 _01000_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[10\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11220_ _03938_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__clkbuf_4
X_20418_ net136 _00449_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[7\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_153_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21398_ net83 _01414_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11151_ _03834_ _03869_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__or2_1
XFILLER_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20349_ rbzero.wall_tracer.rayAddendY\[-7\] _03260_ _09267_ _03276_ vssd1 vssd1 vccd1
+ vccd1 _01416_ sky130_fd_sc_hd__a22o_1
XTAP_6101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11082_ _03782_ _03804_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__and2_1
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14910_ rbzero.wall_tracer.visualWallDist\[2\] _03796_ vssd1 vssd1 vccd1 vccd1 _07524_
+ sky130_fd_sc_hd__nand2_2
XFILLER_118_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15890_ _07861_ _07866_ vssd1 vssd1 vccd1 vccd1 _08504_ sky130_fd_sc_hd__or2b_1
XTAP_5455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ _03795_ rbzero.wall_tracer.stepDistY\[1\] _07450_ _07454_ _04928_ vssd1 vssd1
+ vccd1 vccd1 _07455_ sky130_fd_sc_hd__o221ai_4
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17560_ _10094_ _10096_ vssd1 vssd1 vccd1 vccd1 _10097_ sky130_fd_sc_hd__nand2_1
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14772_ _04927_ rbzero.wall_tracer.stepDistX\[-5\] vssd1 vssd1 vccd1 vccd1 _07386_
+ sky130_fd_sc_hd__nor2_1
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11984_ net16 net15 vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__nor2_1
XFILLER_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16511_ _09118_ _09119_ vssd1 vssd1 vccd1 vccd1 _09120_ sky130_fd_sc_hd__nor2_1
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13723_ _06266_ _06331_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__or2_1
X_17491_ _09345_ _09898_ _09899_ _09274_ _10028_ vssd1 vssd1 vccd1 vccd1 _10029_ sky130_fd_sc_hd__o311a_1
XFILLER_189_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10935_ rbzero.tex_b0\[31\] rbzero.tex_b0\[30\] _03693_ vssd1 vssd1 vccd1 vccd1 _03695_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19230_ _02797_ vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__clkbuf_1
X_16442_ _08398_ _09051_ vssd1 vssd1 vccd1 vccd1 _09052_ sky130_fd_sc_hd__nor2_1
XFILLER_232_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13654_ _06342_ vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__clkbuf_4
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10866_ _03658_ vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ _03816_ _05069_ _05112_ _05293_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__a31o_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19161_ rbzero.spi_registers.new_sky\[1\] rbzero.color_sky\[1\] _02752_ vssd1 vssd1
+ vccd1 vccd1 _02755_ sky130_fd_sc_hd__mux2_1
XFILLER_223_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16373_ _07515_ _08723_ vssd1 vssd1 vccd1 vccd1 _08983_ sky130_fd_sc_hd__nor2_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13585_ _06234_ _06272_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__or2_1
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10797_ _03622_ vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__clkbuf_1
X_18112_ _01796_ _01758_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__or2b_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15324_ _07935_ _07937_ vssd1 vssd1 vccd1 vccd1 _07938_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12536_ _05155_ _05158_ _05156_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__o21a_1
X_19092_ rbzero.spi_registers.mosi rbzero.spi_registers.mosi_buffer\[0\] _04920_ vssd1
+ vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__mux2_1
XFILLER_157_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18043_ rbzero.wall_tracer.trackDistX\[9\] rbzero.wall_tracer.stepDistX\[9\] vssd1
+ vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__nand2_1
X_15255_ _07856_ _07857_ _07868_ vssd1 vssd1 vccd1 vccd1 _07869_ sky130_fd_sc_hd__nand3_1
X_12467_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__nand2_1
XFILLER_126_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14206_ _06862_ _06888_ vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__nand2_1
X_11418_ rbzero.tex_r1\[45\] rbzero.tex_r1\[44\] _03936_ vssd1 vssd1 vccd1 vccd1 _04136_
+ sky130_fd_sc_hd__mux2_1
X_15186_ _07550_ vssd1 vssd1 vccd1 vccd1 _07800_ sky130_fd_sc_hd__buf_2
XFILLER_193_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12398_ _05074_ _05090_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__and2_1
XFILLER_126_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14137_ _06310_ _06634_ vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__nor2_1
XFILLER_119_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11349_ rbzero.row_render.size\[9\] _04048_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__nand2_1
XFILLER_158_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19994_ _03122_ vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__clkinv_2
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14068_ _06741_ _06747_ vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__xor2_1
X_18945_ rbzero.pov.spi_buffer\[21\] rbzero.pov.ready_buffer\[21\] _02629_ vssd1 vssd1
+ vccd1 vccd1 _02632_ sky130_fd_sc_hd__mux2_1
XFILLER_84_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13019_ _05706_ _05707_ _05625_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__a21oi_1
X_18876_ _02576_ _02587_ _02589_ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a21boi_1
XFILLER_95_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17827_ _01498_ _01504_ _01609_ vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__a21oi_1
XFILLER_227_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17758_ _01539_ _01541_ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__or2_1
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16709_ _09257_ vssd1 vssd1 vccd1 vccd1 _09267_ sky130_fd_sc_hd__buf_4
X_17689_ _09182_ _09978_ _01472_ _01473_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__or4bb_1
XFILLER_165_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19428_ _02880_ vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_222_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19359_ _02858_ vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__clkinv_2
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21321_ _00344_ _01337_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21252_ _00301_ _01268_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20203_ _03216_ _03217_ _03218_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__o21ai_1
XFILLER_117_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21183_ _00232_ _01199_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20134_ _03163_ _03164_ _03165_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__or3_1
XFILLER_172_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20065_ _03129_ vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__clkinv_2
XFILLER_86_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20967_ net91 _00983_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ rbzero.tex_g1\[4\] rbzero.tex_g1\[5\] _03574_ vssd1 vssd1 vccd1 vccd1 _03582_
+ sky130_fd_sc_hd__mux2_1
XFILLER_207_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20898_ net60 _00914_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10651_ rbzero.tex_g1\[37\] rbzero.tex_g1\[38\] _03541_ vssd1 vssd1 vccd1 vccd1 _03546_
+ sky130_fd_sc_hd__mux2_1
XFILLER_224_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13370_ _06037_ _06057_ _06058_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__a21oi_1
X_10582_ _03509_ vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12321_ _05008_ _05014_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__nor2_1
XFILLER_155_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15040_ _07647_ _07653_ vssd1 vssd1 vccd1 vccd1 _07654_ sky130_fd_sc_hd__xnor2_1
X_12252_ rbzero.wall_tracer.trackDistX\[1\] _04944_ _04945_ rbzero.wall_tracer.trackDistX\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__o22a_1
XFILLER_177_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11203_ _03911_ _03917_ _03921_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__mux2_1
X_12183_ net36 net37 _04872_ net38 _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__o221a_1
XFILLER_155_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11134_ _03848_ _03851_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__xnor2_1
X_16991_ _07516_ _09114_ vssd1 vssd1 vccd1 vccd1 _09532_ sky130_fd_sc_hd__nor2_1
XFILLER_155_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15942_ _07637_ _07925_ _07924_ vssd1 vssd1 vccd1 vccd1 _08556_ sky130_fd_sc_hd__o21ba_1
XFILLER_153_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11065_ _03789_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__clkbuf_4
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18730_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__nand2_1
XTAP_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18661_ _02390_ _02391_ _02157_ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__a21oi_1
X_15873_ _07840_ _08335_ _08485_ _07838_ vssd1 vssd1 vccd1 vccd1 _08487_ sky130_fd_sc_hd__a2bb2o_1
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17612_ _09345_ _10033_ _10034_ _09274_ _10148_ vssd1 vssd1 vccd1 vccd1 _10149_ sky130_fd_sc_hd__o311a_1
X_14824_ _07336_ _07437_ vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__nand2_1
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18592_ _02330_ _02331_ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__and2_1
XFILLER_224_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17543_ _10071_ _10079_ vssd1 vssd1 vccd1 vccd1 _10080_ sky130_fd_sc_hd__xnor2_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14755_ rbzero.wall_tracer.rayAddendX\[-4\] rbzero.wall_tracer.rayAddendX\[-3\] rbzero.wall_tracer.rayAddendX\[-2\]
+ _05258_ vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__or4_1
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ net18 vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__inv_2
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13706_ _06374_ _06394_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__nor2_1
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17474_ _09874_ _09876_ vssd1 vssd1 vccd1 vccd1 _10012_ sky130_fd_sc_hd__nor2_1
XFILLER_220_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10918_ rbzero.tex_b0\[39\] rbzero.tex_b0\[38\] _03682_ vssd1 vssd1 vccd1 vccd1 _03686_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14686_ _07317_ vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11898_ _04610_ vssd1 vssd1 vccd1 vccd1 o_tex_out0 sky130_fd_sc_hd__buf_2
X_16425_ _08907_ _08908_ _08906_ vssd1 vssd1 vccd1 vccd1 _09035_ sky130_fd_sc_hd__a21o_1
XFILLER_220_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19213_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.new_sky\[1\] _02786_
+ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__mux2_1
XFILLER_204_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13637_ _06325_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__dlymetal6s2s_1
X_10849_ rbzero.tex_g0\[8\] rbzero.tex_g0\[7\] _03649_ vssd1 vssd1 vccd1 vccd1 _03650_
+ sky130_fd_sc_hd__mux2_1
XFILLER_242_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19144_ rbzero.spi_registers.got_new_leak _02724_ vssd1 vssd1 vccd1 vccd1 _02745_
+ sky130_fd_sc_hd__nand2_1
X_16356_ rbzero.wall_tracer.texu\[3\] _07338_ _07266_ _08966_ vssd1 vssd1 vccd1 vccd1
+ _00484_ sky130_fd_sc_hd__o211a_1
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13568_ _06225_ _06255_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__nor2_1
XFILLER_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15307_ _07919_ _07920_ vssd1 vssd1 vccd1 vccd1 _07921_ sky130_fd_sc_hd__or2_1
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12519_ _05155_ _05158_ _05206_ _05207_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__o31a_2
XFILLER_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19075_ rbzero.spi_registers.spi_buffer\[9\] rbzero.spi_registers.spi_buffer\[8\]
+ _02690_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__mux2_1
X_16287_ _08896_ _08897_ vssd1 vssd1 vccd1 vccd1 _08898_ sky130_fd_sc_hd__xnor2_2
XFILLER_173_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13499_ _05621_ _05610_ _06185_ _06186_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__o22a_1
XFILLER_51_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18026_ _01802_ _01803_ _01807_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__a21oi_1
XFILLER_172_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15238_ _07830_ _07850_ _07851_ vssd1 vssd1 vccd1 vccd1 _07852_ sky130_fd_sc_hd__nand3_1
XFILLER_12_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ _07756_ _07781_ vssd1 vssd1 vccd1 vccd1 _07783_ sky130_fd_sc_hd__xor2_1
XFILLER_160_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19977_ _03120_ vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__clkinv_2
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18928_ rbzero.pov.spi_buffer\[13\] rbzero.pov.ready_buffer\[13\] _02618_ vssd1 vssd1
+ vccd1 vccd1 _02623_ sky130_fd_sc_hd__mux2_1
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18859_ _03730_ _02574_ _02568_ vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__o21ai_1
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20821_ _00039_ _00837_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20752_ net105 _00768_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20683_ net76 _00699_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21304_ net128 _01320_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21235_ _00284_ _01251_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21166_ _00215_ _01182_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20117_ _03150_ _03151_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__xnor2_1
XFILLER_132_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21097_ _00146_ _01113_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_219_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20048_ _03125_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__buf_4
XFILLER_213_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12870_ _05406_ _05514_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__nor2_1
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11821_ _03898_ _04526_ _04534_ _03953_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__o211a_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _07099_ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__buf_4
XFILLER_148_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _04323_ _04464_ _04465_ _04466_ _03921_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__o221a_1
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10703_ rbzero.tex_g1\[12\] rbzero.tex_g1\[13\] _03563_ vssd1 vssd1 vccd1 vccd1 _03573_
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14471_ _07102_ _07156_ vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__nand2_1
XFILLER_109_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _03958_ _04396_ _04397_ _04398_ _04007_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__o221a_1
XFILLER_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16210_ _08819_ _08821_ vssd1 vssd1 vccd1 vccd1 _08822_ sky130_fd_sc_hd__xnor2_1
XFILLER_224_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13422_ _06106_ _06110_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__nand2_1
X_17190_ _09467_ _09603_ _09728_ _09729_ vssd1 vssd1 vccd1 vccd1 _09730_ sky130_fd_sc_hd__o31a_1
XFILLER_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10634_ rbzero.tex_g1\[45\] rbzero.tex_g1\[46\] _03530_ vssd1 vssd1 vccd1 vccd1 _03537_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16141_ _08596_ _07886_ vssd1 vssd1 vccd1 vccd1 _08753_ sky130_fd_sc_hd__nor2_1
XFILLER_195_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13353_ _05537_ _05793_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__or2_1
X_10565_ _03500_ vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ rbzero.wall_tracer.trackDistX\[10\] _04995_ rbzero.wall_tracer.trackDistX\[9\]
+ _04991_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__a22o_1
X_16072_ _08659_ _08684_ vssd1 vssd1 vccd1 vccd1 _08685_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13284_ _05971_ _05952_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__and2b_1
XFILLER_108_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10496_ _03464_ vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15023_ _07630_ _07636_ vssd1 vssd1 vccd1 vccd1 _07637_ sky130_fd_sc_hd__nand2_1
XFILLER_182_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19900_ _03112_ vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__clkinv_2
X_12235_ _04930_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__clkbuf_4
XFILLER_216_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19831_ _03106_ vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__clkinv_2
X_12166_ _04871_ net35 vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__nor2_1
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11117_ _03829_ _03835_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__nand2_1
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19762_ _02608_ _03071_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__and2_1
XFILLER_231_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16974_ _09118_ _09500_ vssd1 vssd1 vccd1 vccd1 _09515_ sky130_fd_sc_hd__nand2_1
X_12097_ net43 _04799_ _04802_ _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__a211o_1
XFILLER_96_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18713_ _02434_ _02438_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__nand2_1
XFILLER_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15925_ _07616_ _07914_ vssd1 vssd1 vccd1 vccd1 _08539_ sky130_fd_sc_hd__nor2_1
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11048_ rbzero.otherx\[4\] rbzero.map_rom.i_col\[4\] vssd1 vssd1 vccd1 vccd1 _03776_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_110_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19693_ rbzero.debug_overlay.playerY\[4\] _03043_ vssd1 vssd1 vccd1 vccd1 _03049_
+ sky130_fd_sc_hd__nor2_1
Xinput8 i_gpout0_sel[5] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_4
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15856_ _08468_ _08469_ vssd1 vssd1 vccd1 vccd1 _08470_ sky130_fd_sc_hd__nor2_1
X_18644_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.wall_tracer.rayAddendY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__or2_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14807_ _07351_ rbzero.wall_tracer.stepDistY\[-6\] _07352_ vssd1 vssd1 vccd1 vccd1
+ _07421_ sky130_fd_sc_hd__a21oi_2
XFILLER_40_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15787_ _08399_ _08400_ vssd1 vssd1 vccd1 vccd1 _08401_ sky130_fd_sc_hd__and2_1
X_18575_ _02314_ _02315_ _02305_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__a21oi_1
X_12999_ _05680_ _05682_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__nand2_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17526_ _09797_ _09920_ vssd1 vssd1 vccd1 vccd1 _10063_ sky130_fd_sc_hd__nand2_1
X_14738_ rbzero.wall_tracer.state\[6\] vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__buf_4
XFILLER_205_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17457_ _09985_ _09986_ _09992_ _09993_ vssd1 vssd1 vccd1 vccd1 _09995_ sky130_fd_sc_hd__o22ai_1
XFILLER_127_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14669_ _07308_ vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16408_ _07439_ _07440_ vssd1 vssd1 vccd1 vccd1 _09018_ sky130_fd_sc_hd__nand2_2
XFILLER_242_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17388_ _08890_ _08723_ _09798_ _09799_ vssd1 vssd1 vccd1 vccd1 _09926_ sky130_fd_sc_hd__o31a_1
XFILLER_158_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16339_ _08810_ _08812_ vssd1 vssd1 vccd1 vccd1 _08950_ sky130_fd_sc_hd__nor2_1
XFILLER_186_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19127_ rbzero.othery\[0\] _02723_ _02733_ _02728_ vssd1 vssd1 vccd1 vccd1 _00737_
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19058_ _02691_ vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18009_ _01669_ _01677_ _01790_ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21020_ net94 _01036_ vssd1 vssd1 vccd1 vccd1 rbzero.hsync sky130_fd_sc_hd__dfxtp_1
XFILLER_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20804_ _00022_ _00820_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20735_ net107 _00751_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20666_ net61 _00682_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20597_ net80 _00613_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_109_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10350_ _03385_ vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10281_ _03349_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12020_ net6 _04723_ _04725_ _04728_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__o211a_1
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21218_ _00267_ _01234_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21149_ _00198_ _01165_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_232_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13971_ _06648_ _06654_ vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__and2_1
XFILLER_232_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15710_ _07435_ _08256_ _07592_ _07970_ vssd1 vssd1 vccd1 vccd1 _08324_ sky130_fd_sc_hd__or4_2
X_12922_ _05564_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__buf_2
X_16690_ rbzero.traced_texa\[-6\] _09262_ _09263_ rbzero.wall_tracer.visualWallDist\[-6\]
+ vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__a22o_1
XFILLER_46_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15641_ _08253_ _08254_ vssd1 vssd1 vccd1 vccd1 _08255_ sky130_fd_sc_hd__xor2_1
XFILLER_111_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12853_ _05483_ _05475_ _05478_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__mux2_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ rbzero.wall_tracer.trackDistY\[8\] rbzero.wall_tracer.stepDistY\[8\] vssd1
+ vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__nor2_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11804_ _03825_ _04516_ _04518_ _04117_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__a31o_4
XFILLER_215_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15572_ _08154_ _08156_ vssd1 vssd1 vccd1 vccd1 _08186_ sky130_fd_sc_hd__nor2_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _05462_ _05472_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__nor2_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _09467_ _09603_ _09728_ _09465_ vssd1 vssd1 vccd1 vccd1 _09850_ sky130_fd_sc_hd__o31a_1
XFILLER_15_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14523_ _07200_ vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__clkbuf_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18291_ _02052_ _02054_ _02053_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__a21boi_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11735_ _04448_ _04449_ _03968_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__mux2_1
XFILLER_72_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _09780_ vssd1 vssd1 vccd1 vccd1 _09781_ sky130_fd_sc_hd__inv_2
XFILLER_230_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14454_ _05517_ _07112_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__nand2_1
XFILLER_202_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11666_ _03958_ _04379_ _04380_ _04381_ _04007_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__o221a_1
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13405_ _06089_ _06092_ _06093_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17173_ _09705_ _09712_ vssd1 vssd1 vccd1 vccd1 _09713_ sky130_fd_sc_hd__nand2_1
XFILLER_31_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10617_ rbzero.tex_g1\[53\] rbzero.tex_g1\[54\] _03519_ vssd1 vssd1 vccd1 vccd1 _03528_
+ sky130_fd_sc_hd__mux2_1
X_14385_ _05408_ _07069_ _07073_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__a21oi_1
X_11597_ rbzero.tex_g0\[30\] _04168_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__and2_1
XFILLER_200_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16124_ _07878_ _08735_ vssd1 vssd1 vccd1 vccd1 _08736_ sky130_fd_sc_hd__nor2_1
X_13336_ _06023_ _06024_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__and2_1
XFILLER_182_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10548_ rbzero.tex_r0\[23\] rbzero.tex_r0\[22\] _03490_ vssd1 vssd1 vccd1 vccd1 _03492_
+ sky130_fd_sc_hd__mux2_1
XFILLER_227_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16055_ _07880_ _07620_ rbzero.wall_tracer.visualWallDist\[4\] vssd1 vssd1 vccd1
+ vccd1 _08668_ sky130_fd_sc_hd__or3b_1
XFILLER_143_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13267_ _05912_ _05915_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10479_ _03455_ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__clkbuf_1
X_15006_ _07519_ _07619_ vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__or2_2
X_12218_ _04921_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13198_ _05553_ _05640_ _05651_ _05692_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__a22o_1
XFILLER_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19814_ _02863_ vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__clkinv_2
XFILLER_155_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12149_ net49 net40 net39 net41 _04825_ _04820_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__mux4_1
XFILLER_111_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19745_ rbzero.pov.ready_buffer\[17\] _03067_ _03068_ rbzero.debug_overlay.vplaneX\[-3\]
+ _03015_ vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__a221o_1
X_16957_ _09120_ _09225_ _09498_ vssd1 vssd1 vccd1 vccd1 _09499_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15908_ _08512_ _08521_ vssd1 vssd1 vccd1 vccd1 _08522_ sky130_fd_sc_hd__xor2_2
X_19676_ rbzero.debug_overlay.playerY\[0\] _03016_ _03035_ _03031_ vssd1 vssd1 vccd1
+ vccd1 _00984_ sky130_fd_sc_hd__o211a_1
X_16888_ _09428_ _09429_ _08893_ _09163_ vssd1 vssd1 vccd1 vccd1 _09430_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_225_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18627_ _03737_ _07491_ _02356_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__o21a_1
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15839_ _08172_ _08221_ _08320_ vssd1 vssd1 vccd1 vccd1 _08453_ sky130_fd_sc_hd__and3b_1
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18558_ _02274_ rbzero.wall_tracer.rayAddendX\[7\] vssd1 vssd1 vccd1 vccd1 _02300_
+ sky130_fd_sc_hd__or2_1
XFILLER_75_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17509_ _10044_ _10045_ vssd1 vssd1 vccd1 vccd1 _10046_ sky130_fd_sc_hd__nor2_1
XFILLER_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18489_ _02215_ _02225_ _02210_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__a21bo_1
XANTENNA_13 _07840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20520_ net129 _00536_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_24 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_35 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20451_ net119 _00002_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20382_ net121 _00413_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21003_ net57 _01019_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_5818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11520_ _03783_ _04232_ _04207_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__and3_2
XFILLER_145_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20718_ net93 _00734_ vssd1 vssd1 vccd1 vccd1 rbzero.otherx\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_212_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11451_ rbzero.tex_r1\[29\] rbzero.tex_r1\[28\] _04168_ vssd1 vssd1 vccd1 vccd1 _04169_
+ sky130_fd_sc_hd__mux2_1
X_20649_ net63 _00665_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10402_ _03413_ vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__clkbuf_1
X_14170_ _06470_ _06422_ vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__or2_1
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11382_ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__clkbuf_4
XFILLER_192_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13121_ _05611_ _05607_ _05715_ _05610_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__o22ai_1
XFILLER_152_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10333_ _03376_ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13052_ _05433_ _05740_ _05638_ _05624_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__o22a_1
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10264_ _03340_ vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12003_ net17 _04677_ _04707_ _04712_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__a31o_1
X_17860_ _01635_ _01642_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__xor2_1
XFILLER_117_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10195_ _03304_ vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_105_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16811_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.stepDistX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _09355_ sky130_fd_sc_hd__nor2_1
XFILLER_121_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17791_ _08240_ _09978_ _01460_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__o21bai_1
XFILLER_78_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19530_ rbzero.pov.spi_buffer\[60\] rbzero.pov.spi_buffer\[61\] _02932_ vssd1 vssd1
+ vccd1 vccd1 _02934_ sky130_fd_sc_hd__mux2_1
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13954_ _05740_ _06330_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__nor2_1
X_16742_ _08450_ _08452_ _09293_ _09279_ vssd1 vssd1 vccd1 vccd1 _09294_ sky130_fd_sc_hd__a211oi_4
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12905_ _05314_ _05593_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__nor2_1
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16673_ rbzero.row_render.size\[9\] _09260_ _07206_ _09259_ vssd1 vssd1 vccd1 vccd1
+ _00507_ sky130_fd_sc_hd__a22o_1
XFILLER_62_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19461_ _02897_ vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__clkbuf_1
XFILLER_234_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13885_ _06505_ _06561_ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__xor2_1
XFILLER_235_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18412_ _02163_ _02164_ _02157_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a21oi_1
X_15624_ _08228_ _08230_ vssd1 vssd1 vccd1 vccd1 _08238_ sky130_fd_sc_hd__xor2_1
X_12836_ _05470_ _05514_ _05520_ _05447_ _05524_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__a221oi_4
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19392_ _02861_ vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__clkinv_2
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18343_ _02101_ _02102_ _02103_ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__o21a_1
XFILLER_188_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15555_ _08111_ _08168_ vssd1 vssd1 vccd1 vccd1 _08169_ sky130_fd_sc_hd__nand2_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12767_ _05323_ _05325_ _05448_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__mux2_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14506_ _07177_ _07110_ vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__or2_1
XFILLER_128_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18274_ rbzero.wall_tracer.trackDistY\[-5\] _02039_ _02045_ _09331_ vssd1 vssd1 vccd1
+ vccd1 _00572_ sky130_fd_sc_hd__o22a_1
XFILLER_72_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11718_ rbzero.tex_g1\[39\] rbzero.tex_g1\[38\] _03980_ vssd1 vssd1 vccd1 vccd1 _04434_
+ sky130_fd_sc_hd__mux2_1
XFILLER_202_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15486_ _08097_ _08098_ _08099_ vssd1 vssd1 vccd1 vccd1 _08100_ sky130_fd_sc_hd__a21oi_1
XFILLER_148_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12698_ _05369_ _05372_ _05350_ _05375_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__or4_1
XFILLER_202_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14437_ _07042_ _07040_ vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__and2b_1
X_17225_ _09345_ _09764_ vssd1 vssd1 vccd1 vccd1 _09765_ sky130_fd_sc_hd__and2_1
XFILLER_238_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11649_ rbzero.tex_g0\[34\] _03961_ _03929_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__a21o_1
Xinput11 i_gpout1_sel[2] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_4
XFILLER_204_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput22 i_gpout3_sel[1] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_4
Xinput33 i_gpout5_sel[0] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_4
X_17156_ _09662_ _09695_ vssd1 vssd1 vccd1 vccd1 _09696_ sky130_fd_sc_hd__xnor2_1
Xinput44 i_reg_sclk vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__buf_6
XFILLER_200_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14368_ _07029_ _07053_ _07054_ _07056_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__a31o_1
XFILLER_122_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16107_ _07788_ _07616_ _08718_ _08663_ vssd1 vssd1 vccd1 vccd1 _08719_ sky130_fd_sc_hd__or4_1
X_13319_ _06007_ _05635_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__or2_1
X_17087_ _09489_ _09491_ vssd1 vssd1 vccd1 vccd1 _09628_ sky130_fd_sc_hd__or2b_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14299_ _05432_ _06368_ _06979_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__or3_1
XFILLER_196_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16038_ _08491_ _08493_ vssd1 vssd1 vccd1 vccd1 _08651_ sky130_fd_sc_hd__and2_1
XFILLER_192_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17989_ _09833_ _08725_ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__nor2_1
XFILLER_42_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19728_ rbzero.pov.ready_buffer\[26\] _03061_ _03063_ rbzero.debug_overlay.facingY\[-5\]
+ _03066_ vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__a221o_1
XFILLER_26_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19659_ _07406_ _02958_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__nor2_1
XFILLER_65_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20503_ net133 _00519_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20434_ net131 _00465_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20365_ gpout4.clk_div\[1\] gpout4.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__or2_1
XTAP_7017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20296_ _03258_ vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__clkinv_2
XTAP_6316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10951_ rbzero.tex_b0\[23\] rbzero.tex_b0\[22\] _03693_ vssd1 vssd1 vccd1 vccd1 _03703_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13670_ _06357_ _06358_ _06266_ _06312_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10882_ rbzero.tex_b0\[56\] rbzero.tex_b0\[55\] _03660_ vssd1 vssd1 vccd1 vccd1 _03667_
+ sky130_fd_sc_hd__mux2_1
XFILLER_232_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ _05298_ _05300_ _05307_ _05309_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__and4_1
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15340_ _07951_ _07952_ _07953_ vssd1 vssd1 vccd1 vccd1 _07954_ sky130_fd_sc_hd__a21oi_1
XPHY_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12552_ _05148_ _05151_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__and2b_1
XFILLER_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11503_ _04215_ _04220_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__nor2_1
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15271_ _07878_ _07598_ _07884_ vssd1 vssd1 vccd1 vccd1 _07885_ sky130_fd_sc_hd__or3_1
X_12483_ _05145_ _05144_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__or2b_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17010_ _08223_ _07916_ vssd1 vssd1 vccd1 vccd1 _09551_ sky130_fd_sc_hd__nor2_1
XFILLER_184_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14222_ _06909_ _06910_ vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__nand2_1
XFILLER_138_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11434_ rbzero.tex_r1\[33\] rbzero.tex_r1\[32\] _04148_ vssd1 vssd1 vccd1 vccd1 _04152_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14153_ _06833_ _06832_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__or2b_1
XFILLER_125_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11365_ _04043_ _04083_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__nand2_1
XFILLER_193_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13104_ _05672_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__buf_2
XFILLER_153_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10316_ rbzero.tex_b1\[2\] rbzero.tex_b1\[3\] _03366_ vssd1 vssd1 vccd1 vccd1 _03368_
+ sky130_fd_sc_hd__mux2_1
X_14084_ _06758_ _06759_ _06772_ vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__a21o_1
XFILLER_193_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18961_ _02607_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__clkbuf_4
X_11296_ rbzero.tex_r0\[10\] _04013_ _04014_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__a21o_1
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17912_ _01542_ _01545_ _01694_ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__a21oi_2
X_13035_ _05612_ _05701_ _05717_ _05723_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__a31o_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10247_ _03331_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18892_ rbzero.spi_registers.spi_counter\[5\] rbzero.spi_registers.spi_counter\[4\]
+ rbzero.spi_registers.spi_counter\[3\] _02594_ vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__and4_1
XTAP_6850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17843_ _01578_ _01579_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__nor2_1
XFILLER_117_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10178_ _03290_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__clkbuf_4
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17774_ _01430_ _01437_ _01557_ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__a21oi_1
XFILLER_187_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14986_ rbzero.wall_tracer.rayAddendY\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] _07341_
+ vssd1 vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__mux2_1
XFILLER_208_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19513_ rbzero.pov.spi_buffer\[52\] rbzero.pov.spi_buffer\[53\] _02921_ vssd1 vssd1
+ vccd1 vccd1 _02925_ sky130_fd_sc_hd__mux2_1
XFILLER_75_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16725_ _05121_ vssd1 vssd1 vccd1 vccd1 _09279_ sky130_fd_sc_hd__buf_4
XFILLER_47_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13937_ _06623_ _06625_ vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__or2b_1
XFILLER_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19444_ rbzero.pov.spi_buffer\[19\] rbzero.pov.spi_buffer\[20\] _02888_ vssd1 vssd1
+ vccd1 vccd1 _02889_ sky130_fd_sc_hd__mux2_1
X_13868_ _06507_ _06556_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__xnor2_1
X_16656_ _03810_ vssd1 vssd1 vccd1 vccd1 _09254_ sky130_fd_sc_hd__clkbuf_4
XFILLER_179_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15607_ _08218_ _08220_ vssd1 vssd1 vccd1 vccd1 _08221_ sky130_fd_sc_hd__nor2_2
X_12819_ _05372_ _05378_ _05381_ _05375_ _05428_ _05452_ vssd1 vssd1 vccd1 vccd1 _05508_
+ sky130_fd_sc_hd__mux4_1
XFILLER_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19375_ _02860_ vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__clkinv_2
X_16587_ _09194_ _09195_ vssd1 vssd1 vccd1 vccd1 _09196_ sky130_fd_sc_hd__and2_1
X_13799_ _06426_ _06480_ _06484_ _06487_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_16_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18326_ rbzero.wall_tracer.trackDistY\[3\] rbzero.wall_tracer.stepDistY\[3\] vssd1
+ vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__or2_1
XFILLER_241_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15538_ _08150_ _08151_ vssd1 vssd1 vccd1 vccd1 _08152_ sky130_fd_sc_hd__xor2_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15469_ _07260_ _07408_ _04935_ _07350_ vssd1 vssd1 vccd1 vccd1 _08083_ sky130_fd_sc_hd__or4_1
X_18257_ _02027_ _02028_ _02029_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__a21o_1
X_17208_ _09697_ _09747_ vssd1 vssd1 vccd1 vccd1 _09748_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18188_ _01842_ _01965_ _01967_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__o21a_1
XFILLER_200_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17139_ _09572_ _09574_ _09570_ vssd1 vssd1 vccd1 vccd1 _09679_ sky130_fd_sc_hd__a21bo_1
XFILLER_102_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20150_ _03171_ _03175_ _03172_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__o21ai_1
XFILLER_235_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20081_ _03125_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__buf_4
XFILLER_135_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20983_ net65 _00999_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20417_ net136 _00448_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[6\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_175_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21397_ net86 _01413_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_218_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11150_ _03833_ _03827_ _03829_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__and3_1
X_20348_ _02378_ _03275_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__xnor2_1
XTAP_6102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11081_ gpout0.hpos\[2\] gpout0.hpos\[1\] gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1
+ _03804_ sky130_fd_sc_hd__and3_1
XTAP_6146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20279_ _03256_ vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__clkinv_2
XTAP_6157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ _07337_ _07451_ _07452_ _07453_ vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__a31o_1
XFILLER_188_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ _07351_ rbzero.wall_tracer.stepDistY\[-5\] _07352_ vssd1 vssd1 vccd1 vccd1
+ _07385_ sky130_fd_sc_hd__a21oi_2
XFILLER_112_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11983_ net20 _04692_ _04664_ net17 vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__and4bb_1
XFILLER_229_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16510_ _09010_ _09109_ _09117_ vssd1 vssd1 vccd1 vccd1 _09119_ sky130_fd_sc_hd__and3_1
X_13722_ _05567_ _05748_ _06320_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__and3_1
XFILLER_72_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10934_ _03694_ vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17490_ _10020_ _10025_ _10027_ vssd1 vssd1 vccd1 vccd1 _10028_ sky130_fd_sc_hd__a21o_1
XFILLER_229_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16441_ _08629_ rbzero.wall_tracer.stepDistY\[10\] _07694_ _09050_ vssd1 vssd1 vccd1
+ vccd1 _09051_ sky130_fd_sc_hd__a22oi_4
X_13653_ _06222_ _06341_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__nand2_1
XFILLER_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10865_ net50 rbzero.tex_b0\[63\] _03649_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__mux2_1
XFILLER_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12604_ rbzero.wall_tracer.visualWallDist\[11\] _05190_ vssd1 vssd1 vccd1 vccd1 _05293_
+ sky130_fd_sc_hd__and2_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16372_ _08980_ _08981_ vssd1 vssd1 vccd1 vccd1 _08982_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19160_ rbzero.color_sky\[0\] _02752_ _02754_ vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__a21o_1
X_13584_ _06234_ _06272_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__nand2_1
XFILLER_38_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ rbzero.tex_g0\[33\] rbzero.tex_g0\[32\] _03616_ vssd1 vssd1 vccd1 vccd1 _03622_
+ sky130_fd_sc_hd__mux2_1
XFILLER_223_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _01889_ _01891_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__xor2_1
XFILLER_197_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15323_ _07936_ _07718_ vssd1 vssd1 vccd1 vccd1 _07937_ sky130_fd_sc_hd__nor2_1
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ _05220_ _05221_ _05223_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__o21a_1
XFILLER_129_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19091_ _02709_ vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18042_ rbzero.wall_tracer.trackDistX\[9\] rbzero.wall_tracer.stepDistX\[9\] vssd1
+ vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__or2_1
X_15254_ _07859_ _07867_ vssd1 vssd1 vccd1 vccd1 _07868_ sky130_fd_sc_hd__xor2_1
XFILLER_149_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12466_ _05147_ _05148_ _05153_ _05154_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__o31a_2
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14205_ _06882_ _06893_ vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11417_ _03899_ _04126_ _04134_ _03954_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__o211a_1
X_15185_ _07387_ _07424_ _07552_ _07550_ vssd1 vssd1 vccd1 vccd1 _07799_ sky130_fd_sc_hd__or4_1
XFILLER_67_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12397_ _05044_ _05043_ _05047_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__a21o_1
XFILLER_193_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14136_ _06814_ _06824_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__nor2_1
XFILLER_181_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11348_ _03293_ _04050_ _04051_ gpout0.hpos\[9\] _04066_ vssd1 vssd1 vccd1 vccd1
+ _04067_ sky130_fd_sc_hd__a221o_1
XFILLER_10_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19993_ _03122_ vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__clkinv_2
XFILLER_235_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14067_ _06727_ _06726_ _06712_ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__a21o_1
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18944_ _02631_ vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_234_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11279_ _03995_ _03996_ _03997_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__mux2_1
XFILLER_80_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13018_ _05645_ _05567_ _05604_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__a21bo_1
XFILLER_100_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18875_ rbzero.spi_registers.spi_counter\[0\] _02576_ _02588_ _02589_ vssd1 vssd1
+ vccd1 vccd1 _00629_ sky130_fd_sc_hd__o211a_1
XTAP_6680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17826_ _01498_ _01504_ _01609_ vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__and3_1
XFILLER_230_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17757_ _09166_ _08724_ _10171_ _01540_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__o31a_1
XFILLER_130_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14969_ _07581_ _07582_ _07578_ vssd1 vssd1 vccd1 vccd1 _07583_ sky130_fd_sc_hd__o21a_1
XFILLER_235_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16708_ rbzero.traced_texa\[9\] _09266_ _09265_ rbzero.wall_tracer.visualWallDist\[9\]
+ vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__a22o_1
X_17688_ _08272_ _09449_ _09976_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__a21oi_1
XFILLER_169_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19427_ rbzero.pov.spi_buffer\[11\] rbzero.pov.spi_buffer\[12\] _02877_ vssd1 vssd1
+ vccd1 vccd1 _02880_ sky130_fd_sc_hd__mux2_1
X_16639_ _04593_ _04087_ _09245_ vssd1 vssd1 vccd1 vccd1 _09246_ sky130_fd_sc_hd__and3_1
XFILLER_241_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19358_ _02858_ vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__clkinv_2
XFILLER_52_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18309_ rbzero.wall_tracer.trackDistY\[1\] rbzero.wall_tracer.stepDistY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__or2_1
XFILLER_200_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19289_ _02829_ vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21320_ _00343_ _01336_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21251_ _00300_ _01267_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20202_ _03221_ _03222_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__nand2_1
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21182_ _00231_ _01198_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20133_ _03158_ _03160_ _03159_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__a21boi_1
XFILLER_132_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20064_ _03129_ vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__clkinv_2
XFILLER_58_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20966_ net116 _00982_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_54_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20897_ net60 _00913_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10650_ _03545_ vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10581_ rbzero.tex_r0\[7\] rbzero.tex_r0\[6\] _03501_ vssd1 vssd1 vccd1 vccd1 _03509_
+ sky130_fd_sc_hd__mux2_1
XFILLER_220_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12320_ _04998_ _05013_ _04996_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__o21a_1
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12251_ rbzero.wall_tracer.trackDistY\[0\] vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__inv_2
XFILLER_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11202_ _03920_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__buf_4
XFILLER_194_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12182_ net36 net37 _04872_ net38 _04887_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__a221oi_1
XFILLER_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11133_ _03848_ _03851_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__nor2_1
XFILLER_122_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16990_ _09529_ _09530_ vssd1 vssd1 vccd1 vccd1 _09531_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15941_ _08553_ _08554_ vssd1 vssd1 vccd1 vccd1 _08555_ sky130_fd_sc_hd__xnor2_1
XTAP_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11064_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18660_ _02386_ _02387_ _02389_ vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__o21ai_1
XFILLER_209_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15872_ _07646_ _07840_ _08335_ _08485_ vssd1 vssd1 vccd1 vccd1 _08486_ sky130_fd_sc_hd__or4b_1
XTAP_5275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17611_ _03797_ _10146_ _10147_ vssd1 vssd1 vccd1 vccd1 _10148_ sky130_fd_sc_hd__or3b_2
XFILLER_218_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14823_ _05084_ _05221_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__mux2_1
XFILLER_40_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18591_ _02329_ _02325_ _02326_ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__or3_1
XFILLER_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17542_ _10072_ _10078_ vssd1 vssd1 vccd1 vccd1 _10079_ sky130_fd_sc_hd__xnor2_1
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14754_ _05273_ vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__inv_2
X_11966_ net18 _04675_ _04664_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__o21ba_1
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13705_ _06383_ _06384_ _06385_ _06393_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__o22a_1
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10917_ _03685_ vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17473_ _09912_ _10010_ vssd1 vssd1 vccd1 vccd1 _10011_ sky130_fd_sc_hd__xnor2_2
X_14685_ rbzero.wall_tracer.stepDistX\[-3\] _07192_ _07316_ vssd1 vssd1 vccd1 vccd1
+ _07317_ sky130_fd_sc_hd__mux2_1
XFILLER_229_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11897_ o_tex_oeb0 _04602_ _04606_ _04609_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__and4b_4
XFILLER_232_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19212_ _02787_ vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16424_ _09015_ _09033_ vssd1 vssd1 vccd1 vccd1 _09034_ sky130_fd_sc_hd__xnor2_1
X_13636_ _06115_ _06305_ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__and2_1
XFILLER_32_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10848_ _03604_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__clkbuf_4
XFILLER_160_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19143_ _02743_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__clkbuf_2
X_13567_ _06225_ _06255_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__and2_1
XFILLER_158_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16355_ _04933_ _08964_ _08965_ vssd1 vssd1 vccd1 vccd1 _08966_ sky130_fd_sc_hd__or3_1
X_10779_ rbzero.tex_g0\[41\] rbzero.tex_g0\[40\] _03605_ vssd1 vssd1 vccd1 vccd1 _03613_
+ sky130_fd_sc_hd__mux2_1
XFILLER_203_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15306_ _07791_ _07796_ _07918_ vssd1 vssd1 vccd1 vccd1 _07920_ sky130_fd_sc_hd__a21oi_1
XFILLER_158_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12518_ _05169_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__inv_2
XFILLER_34_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16286_ _08760_ _07736_ vssd1 vssd1 vccd1 vccd1 _08897_ sky130_fd_sc_hd__nor2_1
XFILLER_200_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19074_ _02699_ vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__clkbuf_1
X_13498_ _05621_ _05610_ _06185_ _06186_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__nor4_2
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18025_ _01805_ _01806_ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__nand2_1
XFILLER_51_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15237_ _07845_ _07846_ _07849_ vssd1 vssd1 vccd1 vccd1 _07851_ sky130_fd_sc_hd__a21o_1
XFILLER_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12449_ _05127_ _05133_ _05131_ _05122_ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__o211a_1
XFILLER_201_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15168_ _07756_ _07781_ vssd1 vssd1 vccd1 vccd1 _07782_ sky130_fd_sc_hd__nor2_1
XFILLER_172_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14119_ _06746_ _06802_ _06803_ _06807_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__a31oi_1
X_15099_ _07468_ _07712_ vssd1 vssd1 vccd1 vccd1 _07713_ sky130_fd_sc_hd__nor2_1
XFILLER_114_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19976_ _03120_ vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__clkinv_2
XFILLER_140_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18927_ _02622_ vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18858_ rbzero.wall_tracer.rayAddendY\[11\] _02573_ vssd1 vssd1 vccd1 vccd1 _02574_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_68_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17809_ _01590_ _01592_ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__nor2_1
XFILLER_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18789_ rbzero.wall_tracer.rayAddendY\[4\] rbzero.wall_tracer.rayAddendY\[3\] _02510_
+ vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__o21ai_1
XFILLER_227_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20820_ _00038_ _00836_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20751_ net100 _00767_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_done sky130_fd_sc_hd__dfxtp_1
XFILLER_196_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20682_ net75 _00698_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21303_ net127 _01319_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21234_ _00283_ _01250_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21165_ _00214_ _01181_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20116_ _03143_ _03144_ _03145_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__o21ai_1
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21096_ _00145_ _01112_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20047_ _03127_ vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__clkinv_2
XFILLER_246_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _03920_ _04529_ _04533_ _03949_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__a211o_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ rbzero.tex_b0\[47\] _04143_ _04145_ _03916_ vssd1 vssd1 vccd1 vccd1 _04466_
+ sky130_fd_sc_hd__a31o_1
XFILLER_92_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20949_ net116 _00965_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _03572_ vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14470_ _05470_ _07049_ _07155_ vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__a21oi_2
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11682_ rbzero.tex_g1\[7\] _03964_ _03965_ _03997_ vssd1 vssd1 vccd1 vccd1 _04398_
+ sky130_fd_sc_hd__a31o_1
XFILLER_241_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13421_ _06007_ _06108_ _06109_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__a21bo_1
XFILLER_74_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10633_ _03536_ vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16140_ _08749_ _08751_ vssd1 vssd1 vccd1 vccd1 _08752_ sky130_fd_sc_hd__nand2_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13352_ _06006_ _06011_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__xor2_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10564_ rbzero.tex_r0\[15\] rbzero.tex_r0\[14\] _03490_ vssd1 vssd1 vccd1 vccd1 _03500_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12303_ _04993_ _04996_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__nand2_1
X_16071_ _08661_ _08683_ vssd1 vssd1 vccd1 vccd1 _08684_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13283_ _05952_ _05971_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__xnor2_1
XFILLER_202_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10495_ rbzero.tex_r0\[48\] rbzero.tex_r0\[47\] _03457_ vssd1 vssd1 vccd1 vccd1 _03464_
+ sky130_fd_sc_hd__mux2_1
X_15022_ _07622_ _07635_ vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__nor2_1
XFILLER_108_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12234_ o_vsync rbzero.wall_tracer.state\[4\] _03292_ vssd1 vssd1 vccd1 vccd1 _04930_
+ sky130_fd_sc_hd__and3_1
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19830_ _03106_ vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__clkinv_2
XFILLER_64_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12165_ net36 vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__inv_2
XFILLER_68_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11116_ _03827_ _03828_ rbzero.texV\[6\] vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__a21o_1
XFILLER_190_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19761_ _02838_ _02837_ _02843_ rbzero.pov.spi_done vssd1 vssd1 vccd1 vccd1 _03071_
+ sky130_fd_sc_hd__a31o_1
X_16973_ _09497_ _09499_ vssd1 vssd1 vccd1 vccd1 _09514_ sky130_fd_sc_hd__or2_1
X_12096_ net44 _04798_ _04803_ net42 vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__a22o_1
XFILLER_231_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18712_ _02434_ _02438_ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__or2_1
X_15924_ _08535_ _08537_ vssd1 vssd1 vccd1 vccd1 _08538_ sky130_fd_sc_hd__nand2_1
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11047_ _03769_ _03771_ _03772_ _03774_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__and4bb_1
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19692_ _03008_ _03047_ rbzero.debug_overlay.playerY\[4\] vssd1 vssd1 vccd1 vccd1
+ _03048_ sky130_fd_sc_hd__o21ai_1
XFILLER_232_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 i_gpout1_sel[0] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_6
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18643_ rbzero.debug_overlay.vplaneY\[-9\] rbzero.wall_tracer.rayAddendY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__nand2_1
XFILLER_77_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15855_ _08467_ _08462_ vssd1 vssd1 vccd1 vccd1 _08469_ sky130_fd_sc_hd__and2b_1
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14806_ _07417_ _07419_ _07349_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__a21o_1
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18574_ _02274_ rbzero.debug_overlay.vplaneX\[0\] vssd1 vssd1 vccd1 vccd1 _02315_
+ sky130_fd_sc_hd__or2_1
X_15786_ _07880_ _08398_ _08060_ _07826_ vssd1 vssd1 vccd1 vccd1 _08400_ sky130_fd_sc_hd__o22ai_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ _05667_ _05686_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__xor2_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17525_ _10060_ _10061_ vssd1 vssd1 vccd1 vccd1 _10062_ sky130_fd_sc_hd__xor2_1
XFILLER_166_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14737_ rbzero.wall_tracer.state\[13\] vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__clkbuf_4
XFILLER_33_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11949_ o_tex_sclk _04644_ _04658_ _04659_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__a211oi_1
XFILLER_162_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17456_ _09985_ _09986_ _09992_ _09993_ vssd1 vssd1 vccd1 vccd1 _09994_ sky130_fd_sc_hd__or4_1
XFILLER_177_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14668_ rbzero.wall_tracer.stepDistX\[-11\] _07136_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _07308_ sky130_fd_sc_hd__mux2_1
XFILLER_162_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16407_ _08086_ _07591_ _07790_ _07735_ vssd1 vssd1 vccd1 vccd1 _09017_ sky130_fd_sc_hd__or4_1
X_13619_ _05722_ _05818_ _06306_ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__o21a_1
XFILLER_220_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17387_ _09923_ _09924_ vssd1 vssd1 vccd1 vccd1 _09925_ sky130_fd_sc_hd__xnor2_1
XFILLER_242_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14599_ _07245_ _07259_ _07261_ _07251_ vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__o211a_1
XFILLER_146_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19126_ rbzero.spi_registers.new_other\[0\] _02725_ vssd1 vssd1 vccd1 vccd1 _02733_
+ sky130_fd_sc_hd__or2_1
X_16338_ _08881_ _08948_ vssd1 vssd1 vccd1 vccd1 _08949_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19057_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.mosi _02690_ vssd1
+ vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__mux2_1
X_16269_ _08878_ _08879_ vssd1 vssd1 vccd1 vccd1 _08880_ sky130_fd_sc_hd__nand2_1
XFILLER_134_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18008_ _01568_ _01571_ _01676_ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__a21oi_1
XFILLER_156_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19959_ _03114_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__clkbuf_8
XFILLER_87_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20803_ _00021_ _00819_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20734_ net105 _00750_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20665_ net60 _00681_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20596_ net80 _00612_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10280_ rbzero.tex_b1\[19\] rbzero.tex_b1\[20\] _03344_ vssd1 vssd1 vccd1 vccd1 _03349_
+ sky130_fd_sc_hd__mux2_1
XFILLER_219_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21217_ _00266_ _01233_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21148_ _00197_ _01164_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13970_ _06605_ _06617_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__xnor2_1
X_21079_ _00128_ _01095_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12921_ _05609_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__clkbuf_4
XFILLER_246_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15640_ _07260_ _07453_ _07356_ _07481_ vssd1 vssd1 vccd1 vccd1 _08254_ sky130_fd_sc_hd__or4_2
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12852_ _05458_ _05540_ _05459_ _05394_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__o2bb2a_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _04099_ _04517_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__nand2_1
X_15571_ _08183_ _08184_ vssd1 vssd1 vccd1 vccd1 _08185_ sky130_fd_sc_hd__nand2_1
X_12783_ _05394_ _05385_ _05429_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__mux2_1
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17310_ _09593_ _09722_ _09723_ _09724_ vssd1 vssd1 vccd1 vccd1 _09849_ sky130_fd_sc_hd__a2bb2o_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14522_ rbzero.wall_tracer.stepDistY\[-1\] _07199_ _07193_ vssd1 vssd1 vccd1 vccd1
+ _07200_ sky130_fd_sc_hd__mux2_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ rbzero.tex_b0\[61\] rbzero.tex_b0\[60\] _04013_ vssd1 vssd1 vccd1 vccd1 _04449_
+ sky130_fd_sc_hd__mux2_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.stepDistY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__and2_1
XFILLER_15_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _09663_ _09666_ _09664_ vssd1 vssd1 vccd1 vccd1 _09780_ sky130_fd_sc_hd__a21boi_1
XFILLER_109_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14453_ _07107_ _07139_ _05401_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__o21a_1
X_11665_ rbzero.tex_g1\[31\] _03964_ _03965_ _03997_ vssd1 vssd1 vccd1 vccd1 _04381_
+ sky130_fd_sc_hd__a31o_1
XFILLER_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13404_ _06037_ _06057_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__xnor2_1
X_10616_ _03527_ vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__clkbuf_1
X_17172_ _09710_ _09711_ vssd1 vssd1 vccd1 vccd1 _09712_ sky130_fd_sc_hd__xor2_1
XFILLER_186_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14384_ _05408_ _07072_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__nor2_1
XFILLER_168_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11596_ rbzero.tex_g0\[29\] rbzero.tex_g0\[28\] _03935_ vssd1 vssd1 vccd1 vccd1 _04313_
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16123_ _07916_ vssd1 vssd1 vccd1 vccd1 _08735_ sky130_fd_sc_hd__clkbuf_4
X_13335_ _05937_ _05977_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__xor2_1
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10547_ _03491_ vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16054_ _08537_ _08539_ _08535_ vssd1 vssd1 vccd1 vccd1 _08667_ sky130_fd_sc_hd__a21bo_1
X_13266_ _05920_ _05954_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__nor2_1
XFILLER_108_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10478_ rbzero.tex_r0\[56\] rbzero.tex_r0\[55\] _03446_ vssd1 vssd1 vccd1 vccd1 _03455_
+ sky130_fd_sc_hd__mux2_1
X_15005_ rbzero.wall_tracer.visualWallDist\[3\] _03796_ vssd1 vssd1 vccd1 vccd1 _07619_
+ sky130_fd_sc_hd__nand2_4
X_12217_ o_vsync rbzero.wall_tracer.state\[12\] _04920_ vssd1 vssd1 vccd1 vccd1 _04921_
+ sky130_fd_sc_hd__and3_1
XFILLER_170_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13197_ _05626_ _05630_ _05616_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__a21oi_1
XFILLER_194_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19813_ _02863_ vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__clkinv_2
X_12148_ net43 _04849_ _04852_ _04854_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__a211o_1
XFILLER_2_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19744_ rbzero.pov.ready_buffer\[16\] _03069_ _03070_ rbzero.debug_overlay.vplaneX\[-4\]
+ _02832_ vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__o221a_1
X_16956_ _09223_ _09224_ vssd1 vssd1 vccd1 vccd1 _09498_ sky130_fd_sc_hd__nor2_1
X_12079_ _03294_ _03295_ gpout0.vpos\[8\] _04110_ net21 _04781_ vssd1 vssd1 vccd1
+ vccd1 _04787_ sky130_fd_sc_hd__mux4_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15907_ _08519_ _08520_ vssd1 vssd1 vccd1 vccd1 _08521_ sky130_fd_sc_hd__and2b_1
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19675_ rbzero.pov.ready_buffer\[53\] _02958_ _03007_ _03034_ vssd1 vssd1 vccd1 vccd1
+ _03035_ sky130_fd_sc_hd__a211o_1
X_16887_ _07709_ vssd1 vssd1 vccd1 vccd1 _09429_ sky130_fd_sc_hd__buf_2
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18626_ rbzero.map_rom.f1 _07491_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15838_ _08221_ _08320_ _08451_ vssd1 vssd1 vccd1 vccd1 _08452_ sky130_fd_sc_hd__a21o_1
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18557_ _02274_ rbzero.wall_tracer.rayAddendX\[7\] vssd1 vssd1 vccd1 vccd1 _02299_
+ sky130_fd_sc_hd__nand2_1
X_15769_ _08356_ _08382_ vssd1 vssd1 vccd1 vccd1 _08383_ sky130_fd_sc_hd__nor2_1
XFILLER_205_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17508_ _09947_ _10039_ _10043_ vssd1 vssd1 vccd1 vccd1 _10045_ sky130_fd_sc_hd__and3_1
XFILLER_209_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18488_ _02218_ _02221_ _02233_ _03729_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__a31o_1
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17439_ _09467_ _09728_ _09976_ _09465_ vssd1 vssd1 vccd1 vccd1 _09977_ sky130_fd_sc_hd__o31ai_1
XANTENNA_14 _09200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_25 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_36 _07172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_47 net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20450_ net118 _00001_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_186_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19109_ _02720_ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__buf_4
XFILLER_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20381_ net116 _00412_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21002_ net57 _01018_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_88_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20717_ net93 _00733_ vssd1 vssd1 vccd1 vccd1 rbzero.otherx\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11450_ _03903_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__buf_4
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20648_ net66 _00664_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ rbzero.tex_r1\[26\] rbzero.tex_r1\[27\] _03411_ vssd1 vssd1 vccd1 vccd1 _03413_
+ sky130_fd_sc_hd__mux2_1
X_11381_ _04028_ _04031_ _04099_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__mux2_1
XFILLER_165_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20579_ net87 _00595_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13120_ _05789_ _05790_ _05788_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__a21oi_1
XFILLER_137_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10332_ rbzero.tex_r1\[58\] rbzero.tex_r1\[59\] _03366_ vssd1 vssd1 vccd1 vccd1 _03376_
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13051_ _05622_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__clkbuf_4
XFILLER_139_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10263_ rbzero.tex_b1\[27\] rbzero.tex_b1\[28\] _03333_ vssd1 vssd1 vccd1 vccd1 _03340_
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12002_ _04666_ _04710_ _04711_ _04682_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__a22o_1
XFILLER_156_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10194_ rbzero.tex_b1\[60\] rbzero.tex_b1\[61\] _03300_ vssd1 vssd1 vccd1 vccd1 _03304_
+ sky130_fd_sc_hd__mux2_1
XFILLER_120_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16810_ _07332_ _09099_ vssd1 vssd1 vccd1 vccd1 _09354_ sky130_fd_sc_hd__and2_1
XFILLER_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17790_ _07553_ _09611_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__nand2_1
XFILLER_232_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16741_ _09292_ _08452_ _08450_ vssd1 vssd1 vccd1 vccd1 _09293_ sky130_fd_sc_hd__a21oi_1
XFILLER_87_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13953_ _06137_ _06331_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__nor2_1
XFILLER_46_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12904_ _05431_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__inv_2
XFILLER_47_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19460_ rbzero.pov.spi_buffer\[27\] rbzero.pov.spi_buffer\[28\] _02888_ vssd1 vssd1
+ vccd1 vccd1 _02897_ sky130_fd_sc_hd__mux2_1
X_16672_ rbzero.row_render.size\[8\] _09260_ _07202_ _09259_ vssd1 vssd1 vccd1 vccd1
+ _00506_ sky130_fd_sc_hd__a22o_1
XFILLER_35_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13884_ _06563_ _06572_ vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__nand2_1
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18411_ _02160_ _02161_ _02162_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__o21ai_1
XFILLER_235_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15623_ _08232_ _08236_ _08235_ vssd1 vssd1 vccd1 vccd1 _08237_ sky130_fd_sc_hd__a21bo_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _05447_ _05523_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__nor2_1
X_19391_ _02861_ vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__clkinv_2
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _02101_ _02102_ _02103_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__nor3_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15554_ _08112_ _08167_ vssd1 vssd1 vccd1 vccd1 _08168_ sky130_fd_sc_hd__and2_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12766_ _05327_ _05422_ _05448_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__mux2_1
XFILLER_128_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14505_ _07186_ vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18273_ _01997_ _02043_ _02044_ _02013_ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__a31o_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _03968_ _04430_ _04431_ _04432_ _03994_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__o221a_1
X_15485_ _08078_ _08096_ vssd1 vssd1 vccd1 vccd1 _08099_ sky130_fd_sc_hd__nor2_1
X_12697_ _05378_ _05381_ _05385_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__or3_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17224_ _09760_ _09763_ vssd1 vssd1 vccd1 vccd1 _09764_ sky130_fd_sc_hd__xnor2_4
XFILLER_204_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14436_ _05459_ _06368_ _06979_ _07123_ _07107_ vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__o32a_1
XFILLER_128_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11648_ rbzero.tex_g0\[35\] _04142_ _04144_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__and3_1
XFILLER_198_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 i_gpout1_sel[3] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_4
Xinput23 i_gpout3_sel[2] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_4
Xinput34 i_gpout5_sel[1] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_4
XFILLER_204_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput45 i_reset_lock_a vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_8
X_17155_ _09677_ _09694_ vssd1 vssd1 vccd1 vccd1 _09695_ sky130_fd_sc_hd__xor2_2
XFILLER_196_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14367_ _05531_ _07055_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__and2_1
X_11579_ rbzero.debug_overlay.playerX\[-9\] _04240_ _04289_ _04296_ vssd1 vssd1 vccd1
+ vccd1 _04297_ sky130_fd_sc_hd__a211o_1
XFILLER_200_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16106_ _08717_ vssd1 vssd1 vccd1 vccd1 _08718_ sky130_fd_sc_hd__buf_2
X_13318_ _05489_ _05612_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__nand2_1
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17086_ _09566_ _09626_ vssd1 vssd1 vccd1 vccd1 _09627_ sky130_fd_sc_hd__xnor2_1
X_14298_ _05586_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__buf_2
XFILLER_170_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16037_ _08639_ _08649_ vssd1 vssd1 vccd1 vccd1 _08650_ sky130_fd_sc_hd__xnor2_2
XFILLER_87_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13249_ _05883_ _05884_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17988_ _01767_ _01768_ _01769_ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19727_ rbzero.pov.ready_buffer\[25\] _03056_ _03059_ rbzero.debug_overlay.facingY\[-6\]
+ _03065_ vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__o221a_1
X_16939_ _09469_ _09480_ vssd1 vssd1 vccd1 vccd1 _09481_ sky130_fd_sc_hd__xnor2_1
XFILLER_211_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19658_ rbzero.debug_overlay.playerY\[-5\] _03016_ _03022_ _02978_ vssd1 vssd1 vccd1
+ vccd1 _00979_ sky130_fd_sc_hd__o211a_1
XFILLER_237_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18609_ rbzero.map_rom.f4 _02345_ _09274_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__mux2_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19589_ _02956_ _02968_ _02969_ _02780_ vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__o211a_1
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20502_ net129 _00518_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20433_ net131 _00464_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20364_ gpout4.clk_div\[1\] gpout4.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__nand2_1
XFILLER_228_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20295_ _03258_ vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__clkinv_2
XTAP_6317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10950_ _03702_ vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10881_ _03666_ vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _05277_ _05289_ _05304_ _05308_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__or4_1
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ _05149_ _05150_ _05152_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__o21a_1
XFILLER_240_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11502_ _03780_ _03806_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15270_ _07881_ _07883_ vssd1 vssd1 vccd1 vccd1 _07884_ sky130_fd_sc_hd__nand2_1
X_12482_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] _05164_
+ _05169_ _05170_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__a221o_1
XFILLER_32_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14221_ _06894_ _06896_ vssd1 vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__or2_1
X_11433_ _04149_ _04150_ _04014_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__mux2_1
XFILLER_193_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14152_ _06795_ _06840_ vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__and2_1
X_11364_ _04041_ _04042_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__or2_1
XFILLER_67_1307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13103_ _05674_ _05675_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__xor2_1
X_10315_ _03367_ vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__clkbuf_1
X_14083_ _06761_ _06770_ _06771_ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__a21o_1
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18960_ _02639_ vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11295_ _03915_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__buf_4
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17911_ _08135_ _09115_ _01530_ _01693_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__o31a_1
X_13034_ _05525_ _05722_ _05716_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__and3_1
X_10246_ rbzero.tex_b1\[35\] rbzero.tex_b1\[36\] _03322_ vssd1 vssd1 vccd1 vccd1 _03331_
+ sky130_fd_sc_hd__mux2_1
XFILLER_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18891_ _02601_ vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__clkbuf_1
XTAP_6840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17842_ _01623_ _01624_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__nor2_1
XTAP_6873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10177_ gpout0.hpos\[7\] vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__clkbuf_4
XFILLER_67_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17773_ _01431_ _01436_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__and2_1
XFILLER_232_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14985_ _07213_ _07117_ _07346_ vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__a21o_1
XFILLER_47_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19512_ _02924_ vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__clkbuf_1
X_16724_ _08445_ _08448_ _09277_ vssd1 vssd1 vccd1 vccd1 _09278_ sky130_fd_sc_hd__o21a_1
XFILLER_207_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13936_ _06585_ _06600_ _06624_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__o21ai_1
XFILLER_130_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19443_ _02865_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__clkbuf_4
X_16655_ _03296_ _04206_ _09253_ vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13867_ _06537_ _06555_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__nor2_1
XFILLER_228_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15606_ _08173_ _08217_ vssd1 vssd1 vccd1 vccd1 _08220_ sky130_fd_sc_hd__and2_1
XFILLER_16_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12818_ _05418_ _05362_ _05505_ _05506_ _05429_ _05444_ vssd1 vssd1 vccd1 vccd1 _05507_
+ sky130_fd_sc_hd__mux4_1
X_19374_ _02860_ vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__clkinv_2
XFILLER_76_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16586_ _09184_ _09193_ vssd1 vssd1 vccd1 vccd1 _09195_ sky130_fd_sc_hd__or2_1
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ _06486_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__clkinv_2
XFILLER_72_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18325_ rbzero.wall_tracer.trackDistY\[3\] rbzero.wall_tracer.stepDistY\[3\] vssd1
+ vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__nand2_1
XFILLER_128_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15537_ _08066_ _08068_ vssd1 vssd1 vccd1 vccd1 _08151_ sky130_fd_sc_hd__xnor2_1
XFILLER_163_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12749_ _05367_ _05368_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__nor2_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18256_ _02027_ _02028_ _02029_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__nand3_1
XFILLER_124_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15468_ _07384_ _07385_ _07386_ _07645_ vssd1 vssd1 vccd1 vccd1 _08082_ sky130_fd_sc_hd__a211o_1
XFILLER_175_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17207_ _09744_ _09746_ vssd1 vssd1 vccd1 vccd1 _09747_ sky130_fd_sc_hd__xor2_1
XFILLER_204_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14419_ _05432_ _06980_ _06988_ vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__a21bo_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18187_ _01637_ _01743_ _01745_ _01844_ _01966_ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__a311o_1
XFILLER_198_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15399_ _08010_ _08011_ _08012_ vssd1 vssd1 vccd1 vccd1 _08013_ sky130_fd_sc_hd__a21oi_2
X_17138_ _09549_ _09551_ _09548_ vssd1 vssd1 vccd1 vccd1 _09678_ sky130_fd_sc_hd__a21bo_1
XFILLER_239_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17069_ _04939_ rbzero.wall_tracer.stepDistX\[10\] vssd1 vssd1 vccd1 vccd1 _09610_
+ sky130_fd_sc_hd__nand2_2
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20080_ _03130_ vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__clkinv_2
XFILLER_48_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20982_ net65 _00998_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20416_ net135 _00447_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_107_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21396_ net86 _01412_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20347_ _02373_ _02379_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__and2b_1
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11080_ _03783_ _03780_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__or2_1
XFILLER_27_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20278_ _03256_ vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__clkinv_2
XFILLER_66_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14770_ _07381_ _07383_ _07349_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__a21o_1
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ _04665_ _04519_ _04691_ net18 net19 vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__o2111a_1
XFILLER_112_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13721_ _06408_ _06409_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__xor2_1
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10933_ rbzero.tex_b0\[32\] rbzero.tex_b0\[31\] _03693_ vssd1 vssd1 vccd1 vccd1 _03694_
+ sky130_fd_sc_hd__mux2_1
XFILLER_217_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16440_ _07240_ _08919_ _09049_ _07338_ vssd1 vssd1 vccd1 vccd1 _09050_ sky130_fd_sc_hd__a211o_1
XFILLER_204_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13652_ _06176_ _06221_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__nand2_1
X_10864_ _03657_ vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12603_ _03790_ _05291_ _05187_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__o21ai_2
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _08429_ _08852_ vssd1 vssd1 vccd1 vccd1 _08981_ sky130_fd_sc_hd__nor2_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13583_ _05606_ _06271_ _06239_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__o21a_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10795_ _03621_ vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18110_ _01756_ _01797_ _01890_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__a21oi_1
XFILLER_197_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15322_ _07730_ _07732_ vssd1 vssd1 vccd1 vccd1 _07936_ sky130_fd_sc_hd__nand2_2
XFILLER_158_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12534_ _03815_ _05075_ _05083_ _05222_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__a31o_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19090_ net43 rbzero.spi_registers.mosi_buffer\[0\] _02708_ vssd1 vssd1 vccd1 vccd1
+ _02709_ sky130_fd_sc_hd__mux2_1
XFILLER_184_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18041_ _01821_ _01822_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__or2_2
XFILLER_185_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15253_ _07861_ _07866_ vssd1 vssd1 vccd1 vccd1 _07867_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12465_ rbzero.debug_overlay.facingX\[-6\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__nand2_1
XFILLER_149_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14204_ _06435_ _06634_ vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__nor2_1
XFILLER_32_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11416_ _03921_ _04129_ _04133_ _03950_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__a211o_1
X_15184_ _07796_ _07797_ vssd1 vssd1 vccd1 vccd1 _07798_ sky130_fd_sc_hd__and2_1
XFILLER_165_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12396_ _05087_ _05088_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__xnor2_2
XFILLER_181_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14135_ _06816_ _06822_ _06823_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__a21oi_1
X_11347_ _03293_ _04050_ _04064_ _04065_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__o22a_1
XFILLER_99_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19992_ _03114_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__buf_4
XFILLER_181_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14066_ _06727_ _06712_ _06726_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__nand3_1
XFILLER_193_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11278_ _03942_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__clkbuf_4
X_18943_ rbzero.pov.spi_buffer\[20\] rbzero.pov.ready_buffer\[20\] _02629_ vssd1 vssd1
+ vccd1 vccd1 _02631_ sky130_fd_sc_hd__mux2_1
XFILLER_140_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13017_ _05567_ _05605_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__nand2_1
X_10229_ _03299_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__clkbuf_4
XFILLER_45_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18874_ rbzero.spi_registers.ss_buffer\[1\] _03442_ vssd1 vssd1 vccd1 vccd1 _02589_
+ sky130_fd_sc_hd__nor2_2
XTAP_6670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17825_ _01607_ _01608_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__or2b_2
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17756_ _10058_ _10170_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__nand2_1
XFILLER_78_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14968_ _07508_ _07567_ vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__or2_1
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16707_ rbzero.traced_texa\[8\] _09266_ _09265_ rbzero.wall_tracer.visualWallDist\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__a22o_1
X_13919_ _06510_ _06586_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17687_ _08272_ _09449_ _09976_ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__or3_2
XFILLER_81_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14899_ rbzero.wall_tracer.rayAddendY\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] rbzero.wall_tracer.side
+ vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__mux2_1
XFILLER_90_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19426_ _02879_ vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16638_ _03442_ _03808_ vssd1 vssd1 vccd1 vccd1 _09245_ sky130_fd_sc_hd__nor2_4
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19357_ _02858_ vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__clkinv_2
XFILLER_241_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16569_ _09162_ _09177_ vssd1 vssd1 vccd1 vccd1 _09178_ sky130_fd_sc_hd__xnor2_1
XFILLER_204_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18308_ _04945_ _02001_ _02074_ vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19288_ rbzero.spi_registers.new_vshift\[3\] rbzero.spi_registers.spi_buffer\[3\]
+ _02825_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__mux2_1
XFILLER_176_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18239_ rbzero.wall_tracer.trackDistY\[-9\] rbzero.wall_tracer.stepDistY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__or2_1
XFILLER_191_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21250_ _00299_ _01266_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20201_ rbzero.traced_texa\[5\] rbzero.texV\[5\] vssd1 vssd1 vccd1 vccd1 _03222_
+ sky130_fd_sc_hd__nand2_1
XFILLER_11_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21181_ _00230_ _01197_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20132_ rbzero.traced_texa\[-6\] rbzero.texV\[-6\] vssd1 vssd1 vccd1 vccd1 _03164_
+ sky130_fd_sc_hd__and2_1
XFILLER_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20063_ _03129_ vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__clkinv_2
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20965_ net76 _00981_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20896_ net60 _00912_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10580_ _03508_ vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12250_ rbzero.wall_tracer.trackDistY\[1\] vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__inv_2
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11201_ _03919_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__clkbuf_4
XFILLER_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ net35 _04882_ _04886_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__a21oi_1
XFILLER_120_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21379_ net127 _01395_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11132_ rbzero.texV\[3\] _03849_ _03850_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__a21boi_1
XFILLER_190_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15940_ _07906_ _07928_ vssd1 vssd1 vccd1 vccd1 _08554_ sky130_fd_sc_hd__and2_1
XTAP_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11063_ _03788_ _03785_ _03297_ vssd1 vssd1 vccd1 vccd1 o_tex_csb sky130_fd_sc_hd__a21bo_2
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15871_ _07661_ _07662_ _08484_ vssd1 vssd1 vccd1 vccd1 _08485_ sky130_fd_sc_hd__a21bo_1
XTAP_5265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ _10035_ _10026_ _10145_ vssd1 vssd1 vccd1 vccd1 _10147_ sky130_fd_sc_hd__a21o_1
XTAP_5287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14822_ _07100_ _07191_ _07336_ vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__a21o_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18590_ _02325_ _02326_ _02329_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__o21ai_1
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ _10076_ _10077_ vssd1 vssd1 vccd1 vccd1 _10078_ sky130_fd_sc_hd__nand2_1
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14753_ _07365_ _07366_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__nand2_1
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ _03294_ _03295_ gpout0.vpos\[8\] _04110_ net15 _04671_ vssd1 vssd1 vccd1
+ vccd1 _04675_ sky130_fd_sc_hd__mux4_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13704_ _06317_ _06386_ _06343_ _06392_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__o31a_1
X_17472_ _10008_ _10009_ vssd1 vssd1 vccd1 vccd1 _10010_ sky130_fd_sc_hd__nor2_1
XFILLER_233_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10916_ rbzero.tex_b0\[40\] rbzero.tex_b0\[39\] _03682_ vssd1 vssd1 vccd1 vccd1 _03685_
+ sky130_fd_sc_hd__mux2_1
X_14684_ _04931_ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__buf_4
XFILLER_225_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11896_ _04591_ _04592_ _04607_ _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a211o_1
XFILLER_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19211_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.new_sky\[0\] _02786_
+ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__mux2_1
X_16423_ _09016_ _09032_ vssd1 vssd1 vccd1 vccd1 _09033_ sky130_fd_sc_hd__xor2_1
XFILLER_232_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13635_ _06310_ _06314_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__or2_1
XFILLER_71_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ _03648_ vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19142_ rbzero.spi_registers.got_new_leak _02721_ vssd1 vssd1 vccd1 vccd1 _02743_
+ sky130_fd_sc_hd__and2_1
X_16354_ _08585_ _08963_ vssd1 vssd1 vccd1 vccd1 _08965_ sky130_fd_sc_hd__nor2_1
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13566_ _06214_ _06254_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__xor2_1
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10778_ _03612_ vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_200_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15305_ _07791_ _07796_ _07918_ vssd1 vssd1 vccd1 vccd1 _07919_ sky130_fd_sc_hd__and3_1
XFILLER_199_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12517_ _05167_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__inv_2
XFILLER_9_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19073_ rbzero.spi_registers.spi_buffer\[8\] rbzero.spi_registers.spi_buffer\[7\]
+ _02690_ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__mux2_1
X_16285_ _08894_ _08895_ vssd1 vssd1 vccd1 vccd1 _08896_ sky130_fd_sc_hd__nor2_1
XFILLER_173_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13497_ _06115_ _05848_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__and2_1
XFILLER_145_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18024_ _01663_ _01666_ _01804_ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__nand3_1
X_15236_ _07845_ _07846_ _07849_ vssd1 vssd1 vccd1 vccd1 _07850_ sky130_fd_sc_hd__nand3_1
XFILLER_173_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12448_ _03732_ _05114_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15167_ _07773_ _07779_ _07780_ vssd1 vssd1 vccd1 vccd1 _07781_ sky130_fd_sc_hd__a21oi_1
XFILLER_141_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12379_ _05065_ _05066_ _05070_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__a21o_1
XFILLER_119_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14118_ _06743_ _06804_ _06806_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__and3_1
XFILLER_236_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15098_ _07711_ vssd1 vssd1 vccd1 vccd1 _07712_ sky130_fd_sc_hd__clkbuf_4
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19975_ _03120_ vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__clkinv_2
XFILLER_99_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14049_ _06435_ _06423_ _06736_ _06737_ vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__o31ai_2
XFILLER_140_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18926_ rbzero.pov.spi_buffer\[12\] rbzero.pov.ready_buffer\[12\] _02618_ vssd1 vssd1
+ vccd1 vccd1 _02622_ sky130_fd_sc_hd__mux2_1
XFILLER_141_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18857_ _03809_ _02572_ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__nor2_1
XFILLER_227_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17808_ _01591_ _01480_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__nor2_1
XFILLER_209_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18788_ _02509_ vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__buf_2
XFILLER_243_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17739_ _01521_ _01522_ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__and2_1
XFILLER_36_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20750_ net109 _00766_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19409_ _02870_ vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__clkbuf_1
X_20681_ net76 _00697_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21302_ net128 _01318_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21233_ _00282_ _01249_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21164_ _00213_ _01180_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_236_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20115_ _03148_ _03149_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__nand2_1
XFILLER_132_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21095_ _00144_ _01111_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20046_ _03127_ vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__clkinv_2
XFILLER_58_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ rbzero.tex_b0\[46\] _03959_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__and2_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20948_ net77 _00964_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10701_ rbzero.tex_g1\[13\] rbzero.tex_g1\[14\] _03563_ vssd1 vssd1 vccd1 vccd1 _03572_
+ sky130_fd_sc_hd__mux2_1
XFILLER_198_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ rbzero.tex_g1\[6\] _04374_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__and2_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20879_ net59 _00895_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13420_ _05525_ _05668_ _06107_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__a21o_1
XFILLER_70_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10632_ rbzero.tex_g1\[46\] rbzero.tex_g1\[47\] _03530_ vssd1 vssd1 vccd1 vccd1 _03536_
+ sky130_fd_sc_hd__mux2_1
XFILLER_179_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13351_ _06033_ _06039_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__xor2_1
X_10563_ _03499_ vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12302_ _04994_ rbzero.wall_tracer.trackDistX\[11\] rbzero.wall_tracer.trackDistX\[10\]
+ _04995_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__o22a_1
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16070_ _08666_ _08682_ vssd1 vssd1 vccd1 vccd1 _08683_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13282_ _05953_ _05969_ _05970_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ _03463_ vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15021_ _07631_ _07596_ _07633_ _07634_ vssd1 vssd1 vccd1 vccd1 _07635_ sky130_fd_sc_hd__o31a_1
X_12233_ _04929_ _03730_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__nor2_1
XFILLER_135_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12164_ _04829_ _04847_ _04869_ _04870_ o_rgb[22] vssd1 vssd1 vccd1 vccd1 o_gpout[4]
+ sky130_fd_sc_hd__o32a_4
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11115_ _03827_ _03829_ _03833_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16972_ _09508_ _09513_ rbzero.wall_tracer.trackDistX\[0\] _09276_ vssd1 vssd1 vccd1
+ vccd1 _00553_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_150_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12095_ _04773_ net21 vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__nor2_1
XFILLER_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19760_ rbzero.pov.ready_buffer\[10\] _03055_ _03058_ _02510_ _02832_ vssd1 vssd1
+ vccd1 vccd1 _01033_ sky130_fd_sc_hd__o221a_1
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15923_ _07792_ _07621_ _08536_ _07521_ vssd1 vssd1 vccd1 vccd1 _08537_ sky130_fd_sc_hd__a2bb2o_1
X_11046_ rbzero.otherx\[0\] _03742_ _03744_ rbzero.othery\[3\] _03773_ vssd1 vssd1
+ vccd1 vccd1 _03774_ sky130_fd_sc_hd__o221a_1
XFILLER_42_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18711_ _02422_ _02437_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__xnor2_1
XFILLER_231_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19691_ _02833_ _03044_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__nor2_1
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18642_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.wall_tracer.rayAddendY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__nand2_1
XFILLER_231_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15854_ _08462_ _08467_ vssd1 vssd1 vccd1 vccd1 _08468_ sky130_fd_sc_hd__and2b_1
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14805_ _07346_ _07418_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__nand2_1
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ _02275_ rbzero.debug_overlay.vplaneX\[0\] vssd1 vssd1 vccd1 vccd1 _02314_
+ sky130_fd_sc_hd__nand2_1
X_15785_ _07826_ _07880_ _08398_ _08060_ vssd1 vssd1 vccd1 vccd1 _08399_ sky130_fd_sc_hd__or4_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12997_ _05677_ _05685_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__or2_1
XFILLER_149_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17524_ _09684_ _08723_ vssd1 vssd1 vccd1 vccd1 _10061_ sky130_fd_sc_hd__nor2_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14736_ _07345_ _07348_ _07349_ vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__a21o_1
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11948_ gpout1.clk_div\[0\] _04611_ _04618_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__and3b_1
XFILLER_166_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17455_ _09989_ _09990_ _09991_ vssd1 vssd1 vccd1 vccd1 _09993_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ _07307_ vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11879_ gpout0.hpos\[1\] vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__clkbuf_4
XFILLER_242_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16406_ _08904_ _08911_ _08910_ vssd1 vssd1 vccd1 vccd1 _09016_ sky130_fd_sc_hd__a21bo_1
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13618_ _05606_ _06306_ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__nor2_1
X_17386_ _09022_ _08723_ vssd1 vssd1 vccd1 vccd1 _09924_ sky130_fd_sc_hd__nor2_1
XFILLER_203_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14598_ _07260_ _03800_ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__nand2_1
XFILLER_242_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19125_ rbzero.otherx\[4\] _02723_ _02732_ _02728_ vssd1 vssd1 vccd1 vccd1 _00736_
+ sky130_fd_sc_hd__o211a_1
X_16337_ _08945_ _08947_ vssd1 vssd1 vccd1 vccd1 _08948_ sky130_fd_sc_hd__xor2_1
X_13549_ _05692_ _05722_ _06199_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__and3_1
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19056_ _02689_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__clkbuf_4
X_16268_ _08764_ _08848_ _08877_ vssd1 vssd1 vccd1 vccd1 _08879_ sky130_fd_sc_hd__nand3_1
XFILLER_199_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18007_ _01780_ _01788_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__xnor2_1
XFILLER_103_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15219_ _04937_ rbzero.wall_tracer.stepDistX\[2\] vssd1 vssd1 vccd1 vccd1 _07833_
+ sky130_fd_sc_hd__and2_1
XFILLER_195_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16199_ _08653_ _08654_ vssd1 vssd1 vccd1 vccd1 _08811_ sky130_fd_sc_hd__nor2_1
XFILLER_12_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19958_ _03118_ vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__clkinv_2
XFILLER_68_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18909_ rbzero.pov.spi_buffer\[4\] rbzero.pov.ready_buffer\[4\] _02608_ vssd1 vssd1
+ vccd1 vccd1 _02613_ sky130_fd_sc_hd__mux2_1
XFILLER_101_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19889_ _03111_ vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__clkinv_2
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20802_ _00020_ _00818_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20733_ net107 _00749_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20664_ net60 _00680_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20595_ net96 _00611_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.i_col\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21216_ _00265_ _01232_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21147_ _00196_ _01163_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21078_ _00127_ _01094_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12920_ _05608_ _05566_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20029_ _03126_ vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__clkinv_2
XFILLER_219_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _05539_ _05502_ _05462_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__mux2_1
XFILLER_41_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ rbzero.color_sky\[4\] rbzero.color_floor\[4\] _04030_ vssd1 vssd1 vccd1 vccd1
+ _04517_ sky130_fd_sc_hd__mux2_1
X_15570_ _08177_ _08178_ vssd1 vssd1 vccd1 vccd1 _08184_ sky130_fd_sc_hd__xor2_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12782_ _05447_ _05461_ _05468_ _05470_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__a211o_2
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14521_ _07101_ _07198_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__nand2_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ rbzero.tex_b0\[63\] rbzero.tex_b0\[62\] _04013_ vssd1 vssd1 vccd1 vccd1 _04448_
+ sky130_fd_sc_hd__mux2_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _09667_ _09676_ _09674_ vssd1 vssd1 vccd1 vccd1 _09779_ sky130_fd_sc_hd__a21o_1
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14452_ _05517_ _07108_ _07138_ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11664_ rbzero.tex_g1\[30\] _04374_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__and2_1
XFILLER_109_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13403_ _06090_ _06091_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__nand2_1
X_17171_ _09170_ _09576_ _09578_ _09579_ vssd1 vssd1 vccd1 vccd1 _09711_ sky130_fd_sc_hd__o22a_1
XFILLER_35_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10615_ rbzero.tex_g1\[54\] rbzero.tex_g1\[55\] _03519_ vssd1 vssd1 vccd1 vccd1 _03527_
+ sky130_fd_sc_hd__mux2_1
X_14383_ _07029_ _07071_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__nand2_1
XFILLER_31_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11595_ _04310_ _04311_ _03942_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__mux2_1
X_16122_ _08731_ _08733_ vssd1 vssd1 vccd1 vccd1 _08734_ sky130_fd_sc_hd__nand2_1
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13334_ _05981_ _06022_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__nor2_1
X_10546_ rbzero.tex_r0\[24\] rbzero.tex_r0\[23\] _03490_ vssd1 vssd1 vccd1 vccd1 _03491_
+ sky130_fd_sc_hd__mux2_1
XFILLER_109_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16053_ _08664_ _08665_ vssd1 vssd1 vccd1 vccd1 _08666_ sky130_fd_sc_hd__nand2_1
XFILLER_183_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13265_ _05889_ _05919_ _05918_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__o21a_1
XFILLER_157_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10477_ _03454_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15004_ _07617_ vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__buf_2
XFILLER_237_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12216_ _03292_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__buf_4
X_13196_ _05822_ _05824_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19812_ _02863_ vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__clkinv_2
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12147_ net44 _04848_ _04853_ net42 vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a22o_1
XFILLER_123_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19743_ rbzero.pov.ready_buffer\[15\] _03069_ _03070_ rbzero.debug_overlay.vplaneX\[-5\]
+ _03065_ vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__o221a_1
X_16955_ _09382_ _09496_ vssd1 vssd1 vccd1 vccd1 _09497_ sky130_fd_sc_hd__xnor2_1
X_12078_ _03288_ gpout0.hpos\[1\] _04631_ _04632_ net21 _04781_ vssd1 vssd1 vccd1
+ vccd1 _04786_ sky130_fd_sc_hd__mux4_1
XFILLER_42_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15906_ _08517_ _08518_ vssd1 vssd1 vccd1 vccd1 _08520_ sky130_fd_sc_hd__nand2_1
X_11029_ _03736_ rbzero.map_rom.a6 vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__xor2_1
X_16886_ _07509_ vssd1 vssd1 vccd1 vccd1 _09428_ sky130_fd_sc_hd__buf_2
X_19674_ _03032_ _03033_ _02835_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__a21oi_1
XFILLER_237_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15837_ _08172_ _08218_ vssd1 vssd1 vccd1 vccd1 _08451_ sky130_fd_sc_hd__xnor2_1
X_18625_ _02359_ vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__clkbuf_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15768_ _08357_ _08381_ vssd1 vssd1 vccd1 vccd1 _08382_ sky130_fd_sc_hd__nor2_1
X_18556_ _02287_ _02289_ _02290_ _02298_ vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__a31o_1
XFILLER_212_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17507_ _09947_ _10039_ _10043_ vssd1 vssd1 vccd1 vccd1 _10044_ sky130_fd_sc_hd__a21oi_1
XFILLER_206_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14719_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _07334_ sky130_fd_sc_hd__inv_2
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18487_ _02218_ _02221_ _02233_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a21oi_1
X_15699_ _08284_ _08311_ vssd1 vssd1 vccd1 vccd1 _08313_ sky130_fd_sc_hd__nor2_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17438_ _04939_ _09200_ _09731_ vssd1 vssd1 vccd1 vccd1 _09976_ sky130_fd_sc_hd__o21a_4
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_15 _09470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_26 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_37 _07838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_48 _02708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17369_ _09903_ _09905_ vssd1 vssd1 vccd1 vccd1 _09907_ sky130_fd_sc_hd__or2_1
XFILLER_220_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19108_ _04111_ _04252_ _04113_ _02719_ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__and4_4
X_20380_ net116 _00411_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19039_ rbzero.pov.spi_buffer\[66\] rbzero.pov.ready_buffer\[66\] _02673_ vssd1 vssd1
+ vccd1 vccd1 _02681_ sky130_fd_sc_hd__mux2_1
XFILLER_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21001_ net81 _01017_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_86_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20716_ net93 _00732_ vssd1 vssd1 vccd1 vccd1 rbzero.otherx\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20647_ net66 _00663_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10400_ _03412_ vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11380_ rbzero.floor_leak\[5\] _03896_ _04036_ _04037_ _04098_ vssd1 vssd1 vccd1
+ vccd1 _04099_ sky130_fd_sc_hd__a221o_4
XFILLER_221_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20578_ net89 _00594_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10331_ _03375_ vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13050_ _05401_ _05738_ _05652_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__and3_1
X_10262_ _03339_ vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12001_ net49 net40 net39 net41 _04664_ net15 vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__mux4_1
XFILLER_152_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10193_ _03303_ vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16740_ _08453_ vssd1 vssd1 vccd1 vccd1 _09292_ sky130_fd_sc_hd__inv_2
XFILLER_120_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13952_ _06583_ _06640_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__nand2_1
XFILLER_247_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12903_ _05535_ _05461_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__nand2_1
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16671_ rbzero.row_render.size\[7\] _09260_ _07199_ _09259_ vssd1 vssd1 vccd1 vccd1
+ _00505_ sky130_fd_sc_hd__a22o_1
XFILLER_59_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13883_ _06504_ _06562_ vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__or2_1
XFILLER_228_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15622_ _08233_ _08234_ _08235_ vssd1 vssd1 vccd1 vccd1 _08236_ sky130_fd_sc_hd__a21boi_1
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18410_ _02160_ _02161_ _02162_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__or3_1
X_12834_ _05521_ _05522_ _05478_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__mux2_1
X_19390_ _02861_ vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__clkinv_2
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _02095_ _02097_ _02096_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__o21ba_1
XFILLER_163_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15553_ _08114_ _08166_ vssd1 vssd1 vccd1 vccd1 _08167_ sky130_fd_sc_hd__nor2_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12765_ _05449_ _05451_ _05453_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__mux2_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14504_ rbzero.wall_tracer.stepDistY\[-5\] _07185_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _07186_ sky130_fd_sc_hd__mux2_1
XFILLER_128_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18272_ _02040_ _02041_ _02042_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__a21o_1
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ rbzero.tex_g1\[41\] _03964_ _03965_ _03932_ vssd1 vssd1 vccd1 vccd1 _04432_
+ sky130_fd_sc_hd__a31o_1
XFILLER_202_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15484_ _08070_ _08056_ vssd1 vssd1 vccd1 vccd1 _08098_ sky130_fd_sc_hd__xnor2_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12696_ _05255_ _05384_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__xor2_1
XFILLER_124_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17223_ _09369_ _09761_ _09762_ vssd1 vssd1 vccd1 vccd1 _09763_ sky130_fd_sc_hd__a21bo_1
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14435_ _07105_ _07120_ _07122_ vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__o21a_1
XFILLER_175_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11647_ rbzero.tex_g0\[33\] rbzero.tex_g0\[32\] _04000_ vssd1 vssd1 vccd1 vccd1 _04364_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput13 i_gpout1_sel[4] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_8
XFILLER_168_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput24 i_gpout3_sel[3] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_8
X_17154_ _09692_ _09693_ vssd1 vssd1 vccd1 vccd1 _09694_ sky130_fd_sc_hd__nor2_1
XFILLER_200_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput35 i_gpout5_sel[2] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_4
X_14366_ _07003_ _07022_ _05586_ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__mux2_1
XFILLER_190_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11578_ _04291_ _04293_ _04295_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__or3_1
Xinput46 i_reset_lock_b vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_8
X_16105_ _08716_ vssd1 vssd1 vccd1 vccd1 _08717_ sky130_fd_sc_hd__buf_2
XFILLER_128_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13317_ _06001_ _06005_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__xor2_1
XFILLER_143_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17085_ _09623_ _09625_ vssd1 vssd1 vccd1 vccd1 _09626_ sky130_fd_sc_hd__xor2_1
XFILLER_157_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10529_ rbzero.tex_r0\[32\] rbzero.tex_r0\[31\] _03479_ vssd1 vssd1 vccd1 vccd1 _03482_
+ sky130_fd_sc_hd__mux2_1
XFILLER_239_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14297_ _05432_ _06980_ _06984_ _06985_ vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__a211o_1
XFILLER_157_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16036_ _08647_ _08648_ vssd1 vssd1 vccd1 vccd1 _08649_ sky130_fd_sc_hd__xor2_1
XFILLER_115_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13248_ _05904_ _05930_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13179_ _05866_ _05867_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__and2_1
XFILLER_135_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17987_ _09955_ _08531_ _08985_ _09829_ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__o22a_1
XFILLER_42_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19726_ rbzero.pov.ready_buffer\[24\] _03056_ _03059_ rbzero.debug_overlay.facingY\[-7\]
+ _03065_ vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__o221a_1
X_16938_ _09477_ _09479_ vssd1 vssd1 vccd1 vccd1 _09480_ sky130_fd_sc_hd__xnor2_1
XFILLER_244_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19657_ rbzero.pov.ready_buffer\[48\] _02836_ _03008_ _03021_ vssd1 vssd1 vccd1 vccd1
+ _03022_ sky130_fd_sc_hd__a211o_1
X_16869_ _09409_ _09410_ vssd1 vssd1 vccd1 vccd1 _09411_ sky130_fd_sc_hd__xnor2_1
XFILLER_246_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18608_ rbzero.debug_overlay.playerX\[0\] _03742_ _03798_ vssd1 vssd1 vccd1 vccd1
+ _02345_ sky130_fd_sc_hd__mux2_1
XFILLER_65_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19588_ _07340_ _02960_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__nand2_1
XFILLER_20_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18539_ _02261_ _02282_ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20501_ net133 _00517_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20432_ net131 _00463_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20363_ gpout4.clk_div\[0\] _03003_ vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__nor2_1
XFILLER_31_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20294_ _04702_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__buf_4
XTAP_6307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10880_ rbzero.tex_b0\[57\] rbzero.tex_b0\[56\] _03660_ vssd1 vssd1 vccd1 vccd1 _03666_
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ _03815_ _05089_ _05238_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__a21o_1
XPHY_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11501_ rbzero.debug_overlay.facingX\[-5\] _04214_ _04218_ rbzero.debug_overlay.facingX\[-8\]
+ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__a22o_1
XFILLER_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12481_ _05159_ _05161_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__and2_1
XFILLER_71_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14220_ _06894_ _06896_ vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__nand2_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11432_ rbzero.tex_r1\[37\] rbzero.tex_r1\[36\] _04148_ vssd1 vssd1 vccd1 vccd1 _04150_
+ sky130_fd_sc_hd__mux2_1
XFILLER_165_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14151_ _06836_ _06838_ _06839_ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__o21ba_1
XFILLER_153_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11363_ _04044_ _04081_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__nand2_1
XFILLER_67_1319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13102_ _05789_ _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__xor2_1
XFILLER_152_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10314_ rbzero.tex_b1\[3\] rbzero.tex_b1\[4\] _03366_ vssd1 vssd1 vccd1 vccd1 _03367_
+ sky130_fd_sc_hd__mux2_1
X_14082_ _06763_ _06769_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__and2_1
X_11294_ _03904_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__buf_4
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17910_ _01528_ _01529_ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__nand2_1
X_13033_ _05710_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__clkbuf_2
XFILLER_238_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10245_ _03330_ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18890_ _02590_ _02600_ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__and2_1
XTAP_6830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17841_ _01619_ _01622_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__nor2_1
X_10176_ _03288_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__clkbuf_2
XTAP_6874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17772_ _01548_ _01555_ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__xnor2_1
X_14984_ _07597_ vssd1 vssd1 vccd1 vccd1 _07598_ sky130_fd_sc_hd__buf_2
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19511_ rbzero.pov.spi_buffer\[51\] rbzero.pov.spi_buffer\[52\] _02921_ vssd1 vssd1
+ vccd1 vccd1 _02924_ sky130_fd_sc_hd__mux2_1
X_13935_ _06583_ _06601_ vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__or2b_1
X_16723_ _08445_ _08448_ _05121_ vssd1 vssd1 vccd1 vccd1 _09277_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16654_ _03296_ _04206_ _09245_ vssd1 vssd1 vccd1 vccd1 _09253_ sky130_fd_sc_hd__o21ai_1
XFILLER_47_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19442_ _02887_ vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__clkbuf_1
XFILLER_234_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13866_ _06553_ _06554_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__and2b_1
XFILLER_222_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15605_ _08172_ _08218_ vssd1 vssd1 vccd1 vccd1 _08219_ sky130_fd_sc_hd__and2b_1
X_12817_ _05417_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__inv_2
X_16585_ _09184_ _09193_ vssd1 vssd1 vccd1 vccd1 _09194_ sky130_fd_sc_hd__nand2_1
XFILLER_234_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19373_ _02860_ vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__clkinv_2
XFILLER_90_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13797_ _06426_ _06480_ _06485_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18324_ rbzero.wall_tracer.trackDistY\[2\] _02039_ _02088_ _09765_ vssd1 vssd1 vccd1
+ vccd1 _00579_ sky130_fd_sc_hd__o22a_1
X_15536_ _08121_ _08129_ _08149_ vssd1 vssd1 vccd1 vccd1 _08150_ sky130_fd_sc_hd__a21o_1
X_12748_ _05321_ _05383_ _05388_ _05436_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__a31oi_2
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18255_ _02021_ _02023_ _02022_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__o21bai_1
XFILLER_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15467_ _08010_ _08011_ vssd1 vssd1 vccd1 vccd1 _08081_ sky130_fd_sc_hd__xnor2_1
XFILLER_198_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12679_ _05296_ _05263_ _05233_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__a21oi_1
XFILLER_129_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17206_ _09589_ _09622_ _09745_ vssd1 vssd1 vccd1 vccd1 _09746_ sky130_fd_sc_hd__a21boi_1
X_14418_ _05499_ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__buf_2
XFILLER_147_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18186_ _09968_ _01743_ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__and2_1
X_15398_ _08008_ _08009_ vssd1 vssd1 vccd1 vccd1 _08012_ sky130_fd_sc_hd__and2b_1
XFILLER_190_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17137_ _09667_ _09676_ vssd1 vssd1 vccd1 vccd1 _09677_ sky130_fd_sc_hd__xor2_2
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14349_ _07029_ _06987_ _07031_ _07037_ vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__a31o_1
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17068_ _09474_ _09475_ _09201_ vssd1 vssd1 vccd1 vccd1 _09609_ sky130_fd_sc_hd__a21o_1
XFILLER_171_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16019_ _07228_ _08630_ _08631_ _07337_ vssd1 vssd1 vccd1 vccd1 _08632_ sky130_fd_sc_hd__a211o_1
XFILLER_83_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19709_ _02721_ _02954_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__nand2_1
XFILLER_214_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20981_ net90 _00997_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_226_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20415_ net136 _00446_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_175_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21395_ net86 _01411_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20346_ _09257_ _02377_ _03274_ _02158_ rbzero.wall_tracer.rayAddendY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__a32o_1
XFILLER_88_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20277_ _03256_ vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__clkinv_2
XTAP_6126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11981_ _04665_ o_rgb[23] vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__nand2_1
XFILLER_44_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13720_ _06327_ _06378_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10932_ _03604_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__clkbuf_4
XFILLER_84_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13651_ _05767_ _06331_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__nor2_1
XFILLER_147_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10863_ rbzero.tex_g0\[1\] rbzero.tex_g0\[0\] _03649_ vssd1 vssd1 vccd1 vccd1 _03657_
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12602_ _05290_ _03816_ _05188_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__o21a_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16370_ _07625_ _08979_ vssd1 vssd1 vccd1 vccd1 _08980_ sky130_fd_sc_hd__or2_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _06268_ _06270_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ rbzero.tex_g0\[34\] rbzero.tex_g0\[33\] _03616_ vssd1 vssd1 vccd1 vccd1 _03621_
+ sky130_fd_sc_hd__mux2_1
XFILLER_197_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15321_ _07439_ _07440_ _07441_ _07645_ vssd1 vssd1 vccd1 vccd1 _07935_ sky130_fd_sc_hd__a211o_1
XFILLER_158_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12533_ rbzero.wall_tracer.visualWallDist\[-3\] _05189_ rbzero.wall_tracer.rcp_sel\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__a21o_1
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18040_ _01711_ _01720_ _01820_ _03798_ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__a31o_1
XFILLER_184_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15252_ _07864_ _07865_ vssd1 vssd1 vccd1 vccd1 _07866_ sky130_fd_sc_hd__xor2_1
XFILLER_129_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12464_ _05149_ _05150_ _05151_ _05152_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__o211a_1
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14203_ _06858_ _06889_ _06891_ vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__o21ai_1
XFILLER_184_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11415_ _03910_ _04130_ _04131_ _04132_ _03945_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__o221a_1
X_15183_ _07788_ _07598_ _07795_ vssd1 vssd1 vccd1 vccd1 _07797_ sky130_fd_sc_hd__o21ai_1
XFILLER_158_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12395_ _05038_ _05041_ _05042_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__a21o_1
XFILLER_181_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14134_ _06817_ _06821_ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__and2b_1
X_11346_ _03290_ _04052_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__and2_1
XFILLER_180_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19991_ _03121_ vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__clkinv_2
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14065_ _06751_ _06753_ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__nor2_1
X_18942_ _02630_ vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__clkbuf_1
XFILLER_165_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11277_ rbzero.tex_r0\[25\] rbzero.tex_r0\[24\] _03936_ vssd1 vssd1 vccd1 vccd1 _03996_
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13016_ _05703_ _05704_ _05629_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__a21o_1
XFILLER_84_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10228_ _03321_ vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__clkbuf_1
XFILLER_239_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18873_ rbzero.spi_registers.spi_counter\[0\] _02587_ _02576_ vssd1 vssd1 vccd1 vccd1
+ _02588_ sky130_fd_sc_hd__o21ai_1
XTAP_6660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17824_ _01513_ _01514_ _01606_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__a21o_1
XFILLER_227_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17755_ _01537_ _01538_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__xnor2_1
X_14967_ _07578_ _07580_ vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__nand2_1
XFILLER_130_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16706_ _09254_ vssd1 vssd1 vccd1 vccd1 _09266_ sky130_fd_sc_hd__buf_2
X_13918_ _06512_ _06606_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__xor2_1
XFILLER_130_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17686_ _10113_ _10114_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__nand2_1
XFILLER_208_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14898_ _07511_ vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__inv_2
XFILLER_63_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19425_ rbzero.pov.spi_buffer\[10\] rbzero.pov.spi_buffer\[11\] _02877_ vssd1 vssd1
+ vccd1 vccd1 _02879_ sky130_fd_sc_hd__mux2_1
X_13849_ _06484_ _06486_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__xor2_1
X_16637_ _03289_ _09244_ vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__nor2_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19356_ _02858_ vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__clkinv_2
X_16568_ _09168_ _09176_ vssd1 vssd1 vccd1 vccd1 _09177_ sky130_fd_sc_hd__xnor2_1
XFILLER_222_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18307_ _09345_ _02072_ _02073_ _09508_ _01995_ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__o311a_1
XFILLER_52_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15519_ _08122_ _08132_ vssd1 vssd1 vccd1 vccd1 _08133_ sky130_fd_sc_hd__xor2_1
X_16499_ _08968_ _09101_ _09102_ vssd1 vssd1 vccd1 vccd1 _09108_ sky130_fd_sc_hd__a21boi_1
X_19287_ _02828_ vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18238_ rbzero.wall_tracer.trackDistY\[-10\] _01996_ _02014_ _09294_ vssd1 vssd1
+ vccd1 vccd1 _00567_ sky130_fd_sc_hd__o22a_1
XFILLER_136_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18169_ _09833_ _09829_ _08852_ _09373_ vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__or4_1
XFILLER_116_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20200_ rbzero.traced_texa\[5\] rbzero.texV\[5\] vssd1 vssd1 vccd1 vccd1 _03221_
+ sky130_fd_sc_hd__or2_1
XFILLER_85_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21180_ _00229_ _01196_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20131_ rbzero.traced_texa\[-6\] rbzero.texV\[-6\] vssd1 vssd1 vccd1 vccd1 _03163_
+ sky130_fd_sc_hd__nor2_1
XFILLER_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20062_ _03129_ vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__clkinv_2
XFILLER_98_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20964_ net116 _00980_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20895_ net62 _00911_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11200_ _03864_ _03894_ _03918_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__nor3_2
XFILLER_218_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12180_ _04876_ _04884_ _04885_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__o21a_1
X_21378_ net119 _01394_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11131_ rbzero.traced_texVinit\[3\] rbzero.spi_registers.vshift\[0\] vssd1 vssd1
+ vccd1 vccd1 _03850_ sky130_fd_sc_hd__nand2_1
XFILLER_218_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20329_ gpout1.clk_div\[0\] gpout1.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__nand2_1
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11062_ _03290_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__inv_2
XTAP_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15870_ _07466_ rbzero.wall_tracer.stepDistX\[3\] vssd1 vssd1 vccd1 vccd1 _08484_
+ sky130_fd_sc_hd__nand2_1
XTAP_5244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14821_ _07434_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__buf_2
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17540_ _09571_ _08735_ _10075_ vssd1 vssd1 vccd1 vccd1 _10077_ sky130_fd_sc_hd__o21ai_1
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ rbzero.debug_overlay.playerX\[-6\] _07364_ vssd1 vssd1 vccd1 vccd1 _07366_
+ sky130_fd_sc_hd__nand2_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _04591_ _04080_ _04628_ _04101_ _04665_ _04671_ vssd1 vssd1 vccd1 vccd1 _04674_
+ sky130_fd_sc_hd__mux4_1
XFILLER_233_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13703_ _05861_ _06389_ _06391_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__or3b_1
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17471_ _10005_ _10007_ vssd1 vssd1 vccd1 vccd1 _10009_ sky130_fd_sc_hd__and2_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10915_ _03684_ vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__clkbuf_1
X_14683_ _07315_ vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11895_ _03289_ _04604_ _03782_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__a21bo_1
XFILLER_60_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19210_ _02785_ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__clkbuf_4
X_16422_ _09024_ _09031_ vssd1 vssd1 vccd1 vccd1 _09032_ sky130_fd_sc_hd__xnor2_1
X_13634_ _06316_ _06322_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__and2_1
XFILLER_220_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10846_ rbzero.tex_g0\[9\] rbzero.tex_g0\[8\] _03638_ vssd1 vssd1 vccd1 vccd1 _03648_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16353_ _08585_ _08963_ vssd1 vssd1 vccd1 vccd1 _08964_ sky130_fd_sc_hd__and2_1
X_19141_ rbzero.spi_registers.new_vinf _02739_ _02740_ _02741_ _02742_ vssd1 vssd1
+ vccd1 vccd1 _00742_ sky130_fd_sc_hd__o311a_1
XFILLER_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13565_ _06228_ _06253_ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__xnor2_2
XFILLER_201_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10777_ rbzero.tex_g0\[42\] rbzero.tex_g0\[41\] _03605_ vssd1 vssd1 vccd1 vccd1 _03612_
+ sky130_fd_sc_hd__mux2_1
X_15304_ _07913_ _07917_ vssd1 vssd1 vccd1 vccd1 _07918_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12516_ _05159_ _05160_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__nand2_1
X_19072_ _02698_ vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__clkbuf_1
X_16284_ _08240_ _07685_ _07712_ _07800_ vssd1 vssd1 vccd1 vccd1 _08895_ sky130_fd_sc_hd__o22a_1
XFILLER_173_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13496_ _05401_ _06115_ _05848_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18023_ _01663_ _01666_ _01804_ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__a21o_1
XFILLER_195_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15235_ _07663_ _07847_ _07654_ _07848_ vssd1 vssd1 vccd1 vccd1 _07849_ sky130_fd_sc_hd__o31ai_1
X_12447_ _05137_ vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15166_ _07757_ _07772_ vssd1 vssd1 vccd1 vccd1 _07780_ sky130_fd_sc_hd__nor2_1
XFILLER_160_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12378_ _05065_ _05066_ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__and3_1
XFILLER_181_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14117_ _06802_ _06805_ vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11329_ rbzero.row_render.size\[7\] rbzero.row_render.size\[6\] rbzero.row_render.size\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__a21o_1
X_15097_ _07709_ _07710_ vssd1 vssd1 vccd1 vccd1 _07711_ sky130_fd_sc_hd__and2_1
XFILLER_114_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19974_ _03120_ vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__clkinv_2
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14048_ _06734_ _06735_ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__nand2_1
XFILLER_45_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18925_ _02621_ vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18856_ _02570_ _02510_ _02571_ vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__mux2_1
XTAP_6490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17807_ _10120_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__inv_2
XFILLER_227_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18787_ _02472_ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__buf_2
XFILLER_227_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15999_ _08601_ _08611_ vssd1 vssd1 vccd1 vccd1 _08612_ sky130_fd_sc_hd__xor2_2
XFILLER_83_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17738_ _01445_ _01516_ _01520_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__nand3_1
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17669_ _01452_ _01453_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__nand2_1
XFILLER_208_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19408_ rbzero.pov.spi_buffer\[2\] rbzero.pov.spi_buffer\[3\] _02866_ vssd1 vssd1
+ vccd1 vccd1 _02870_ sky130_fd_sc_hd__mux2_1
XFILLER_168_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20680_ net74 _00696_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19339_ _02857_ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__clkinv_2
XFILLER_143_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21301_ net132 _01317_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21232_ _00281_ _01248_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21163_ _00212_ _01179_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20114_ rbzero.traced_texa\[-9\] rbzero.texV\[-9\] vssd1 vssd1 vccd1 vccd1 _03149_
+ sky130_fd_sc_hd__nand2_1
XFILLER_137_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21094_ _00143_ _01110_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20045_ _03127_ vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__clkinv_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ net116 _00963_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10700_ _03571_ vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_230_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ rbzero.tex_g1\[5\] rbzero.tex_g1\[4\] _03962_ vssd1 vssd1 vccd1 vccd1 _04396_
+ sky130_fd_sc_hd__mux2_1
XFILLER_241_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20878_ net58 _00894_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_198_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10631_ _03535_ vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13350_ _06032_ _06034_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__nand2_1
XFILLER_122_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10562_ rbzero.tex_r0\[16\] rbzero.tex_r0\[15\] _03490_ vssd1 vssd1 vccd1 vccd1 _03499_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12301_ rbzero.wall_tracer.trackDistY\[10\] vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__inv_2
XFILLER_127_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13281_ _05968_ _05955_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__and2b_1
X_10493_ rbzero.tex_r0\[49\] rbzero.tex_r0\[48\] _03457_ vssd1 vssd1 vccd1 vccd1 _03463_
+ sky130_fd_sc_hd__mux2_1
X_15020_ _07594_ _07595_ vssd1 vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__nand2_1
XFILLER_68_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12232_ _04928_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__buf_4
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12163_ _04830_ _04853_ _04860_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__nand3_1
XFILLER_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11114_ rbzero.texV\[7\] _03832_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16971_ _07332_ _09511_ _09512_ _09275_ vssd1 vssd1 vccd1 vccd1 _09513_ sky130_fd_sc_hd__o31a_1
X_12094_ _04773_ net21 _04116_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__and3_1
XFILLER_231_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18710_ _02435_ _02436_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__nor2_1
XFILLER_81_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15922_ _04938_ _07617_ vssd1 vssd1 vccd1 vccd1 _08536_ sky130_fd_sc_hd__nor2_2
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11045_ rbzero.othery\[0\] rbzero.map_rom.d6 vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__xnor2_1
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19690_ rbzero.debug_overlay.playerY\[3\] _03008_ _03046_ _02989_ vssd1 vssd1 vccd1
+ vccd1 _00987_ sky130_fd_sc_hd__a211o_1
XFILLER_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18641_ rbzero.debug_overlay.vplaneY\[-7\] rbzero.wall_tracer.rayAddendY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__nor2_1
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15853_ _08465_ _08466_ vssd1 vssd1 vccd1 vccd1 _08467_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14804_ _05089_ _05236_ _07341_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__mux2_1
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18572_ _02287_ _02303_ _02304_ _02313_ vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__a31o_1
X_15784_ _07971_ vssd1 vssd1 vccd1 vccd1 _08398_ sky130_fd_sc_hd__clkbuf_4
X_12996_ _05682_ _05683_ _05684_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__and3_1
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _10057_ _10059_ vssd1 vssd1 vccd1 vccd1 _10060_ sky130_fd_sc_hd__or2b_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14735_ rbzero.wall_tracer.state\[13\] vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__clkbuf_4
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11947_ _04623_ _04653_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__nand2_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ _09989_ _09990_ _09991_ vssd1 vssd1 vccd1 vccd1 _09992_ sky130_fd_sc_hd__and3_1
X_14666_ rbzero.wall_tracer.stepDistX\[-12\] _07118_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _07307_ sky130_fd_sc_hd__mux2_1
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11878_ gpout0.hpos\[2\] vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__buf_2
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16405_ _08892_ _08900_ _09014_ vssd1 vssd1 vccd1 vccd1 _09015_ sky130_fd_sc_hd__a21o_1
X_13617_ _06305_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__buf_2
XFILLER_158_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10829_ _03639_ vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17385_ _09797_ _09920_ _09922_ vssd1 vssd1 vccd1 vccd1 _09923_ sky130_fd_sc_hd__a21oi_1
X_14597_ rbzero.wall_tracer.visualWallDist\[-10\] vssd1 vssd1 vccd1 vccd1 _07260_
+ sky130_fd_sc_hd__clkinv_2
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19124_ rbzero.spi_registers.new_other\[10\] _02725_ vssd1 vssd1 vccd1 vccd1 _02732_
+ sky130_fd_sc_hd__or2_1
X_16336_ _08767_ _08809_ _08946_ vssd1 vssd1 vccd1 vccd1 _08947_ sky130_fd_sc_hd__a21o_1
XFILLER_192_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13548_ _06184_ _06187_ _06188_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__or3_1
XFILLER_242_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16267_ _08764_ _08848_ _08877_ vssd1 vssd1 vccd1 vccd1 _08878_ sky130_fd_sc_hd__a21o_1
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19055_ rbzero.spi_registers.spi_counter\[3\] rbzero.spi_registers.spi_counter\[2\]
+ _02577_ _02576_ _02589_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__o311a_1
X_13479_ _06155_ _06157_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18006_ _01781_ _01787_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__xnor2_1
X_15218_ _07831_ vssd1 vssd1 vccd1 vccd1 _07832_ sky130_fd_sc_hd__inv_2
XFILLER_173_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16198_ _08767_ _08809_ vssd1 vssd1 vccd1 vccd1 _08810_ sky130_fd_sc_hd__xnor2_1
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15149_ _07759_ _07762_ vssd1 vssd1 vccd1 vccd1 _07763_ sky130_fd_sc_hd__and2_1
XFILLER_236_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19957_ _03118_ vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__clkinv_2
XFILLER_84_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18908_ _02612_ vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19888_ _03111_ vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__clkinv_2
XFILLER_68_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18839_ _02510_ rbzero.wall_tracer.rayAddendY\[9\] vssd1 vssd1 vccd1 vccd1 _02557_
+ sky130_fd_sc_hd__xor2_1
XFILLER_95_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20801_ _00019_ _00817_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_222_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20732_ net103 _00748_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20663_ net67 _00679_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20594_ net92 _00610_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f1 sky130_fd_sc_hd__dfxtp_2
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21215_ _00264_ _01231_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21146_ _00195_ _01162_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21077_ _00126_ _01093_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20028_ _03126_ vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__clkinv_2
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12850_ _05381_ _05375_ _05463_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__mux2_1
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _04099_ _04481_ _04515_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__nand3b_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _05469_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__clkbuf_4
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _05602_ _07080_ _07150_ _07177_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__o2bb2a_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11732_ _04447_ vssd1 vssd1 vccd1 vccd1 o_rgb[15] sky130_fd_sc_hd__inv_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14451_ _05497_ _07104_ vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__or2_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11663_ rbzero.tex_g1\[29\] rbzero.tex_g1\[28\] _04378_ vssd1 vssd1 vccd1 vccd1 _04379_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13402_ _06068_ _06088_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__xnor2_1
X_17170_ _09708_ _09709_ vssd1 vssd1 vccd1 vccd1 _09710_ sky130_fd_sc_hd__xor2_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10614_ _03526_ vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__clkbuf_1
X_14382_ _07041_ _07070_ _05586_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__mux2_1
XFILLER_70_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ rbzero.tex_g0\[25\] rbzero.tex_g0\[24\] _03935_ vssd1 vssd1 vccd1 vccd1 _04311_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16121_ _08599_ _08732_ _08536_ _07882_ vssd1 vssd1 vccd1 vccd1 _08733_ sky130_fd_sc_hd__a2bb2o_1
X_13333_ _05992_ _06020_ _06021_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__a21oi_2
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10545_ _03445_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__clkbuf_4
XFILLER_183_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16052_ _07633_ _08663_ _08662_ vssd1 vssd1 vccd1 vccd1 _08665_ sky130_fd_sc_hd__o21ai_1
X_13264_ _05940_ _05945_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10476_ rbzero.tex_r0\[57\] rbzero.tex_r0\[56\] _03446_ vssd1 vssd1 vccd1 vccd1 _03454_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15003_ rbzero.wall_tracer.visualWallDist\[4\] _03796_ vssd1 vssd1 vccd1 vccd1 _07617_
+ sky130_fd_sc_hd__nand2_1
X_12215_ rbzero.hsync vssd1 vssd1 vccd1 vccd1 o_hsync sky130_fd_sc_hd__inv_2
XFILLER_68_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13195_ _05793_ _05728_ _05819_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__or3_2
XFILLER_124_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19811_ _02863_ vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__clkinv_2
X_12146_ _04825_ net27 vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__nor2_1
XFILLER_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19742_ rbzero.pov.ready_buffer\[14\] _03069_ _03070_ rbzero.debug_overlay.vplaneX\[-6\]
+ _03065_ vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__o221a_1
X_16954_ _09493_ _09495_ vssd1 vssd1 vccd1 vccd1 _09496_ sky130_fd_sc_hd__xor2_1
XFILLER_173_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12077_ net24 vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__inv_2
XFILLER_81_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15905_ _08517_ _08518_ vssd1 vssd1 vccd1 vccd1 _08519_ sky130_fd_sc_hd__nor2_1
X_11028_ rbzero.map_rom.d6 rbzero.map_rom.c6 _03739_ _03750_ _03755_ vssd1 vssd1 vccd1
+ vccd1 _03756_ sky130_fd_sc_hd__a311o_1
X_19673_ rbzero.debug_overlay.playerY\[0\] _07498_ vssd1 vssd1 vccd1 vccd1 _03033_
+ sky130_fd_sc_hd__nand2_1
X_16885_ _07591_ _07509_ _07685_ _07709_ vssd1 vssd1 vccd1 vccd1 _09427_ sky130_fd_sc_hd__or4_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18624_ _03736_ _02358_ _09274_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__mux2_1
XFILLER_168_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15836_ _08221_ _08319_ _08322_ _08449_ vssd1 vssd1 vccd1 vccd1 _08450_ sky130_fd_sc_hd__a22o_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18555_ rbzero.wall_tracer.rayAddendX\[6\] _02197_ _02297_ _02157_ vssd1 vssd1 vccd1
+ vccd1 _02298_ sky130_fd_sc_hd__a22o_1
XFILLER_209_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15767_ _08375_ _08379_ _08380_ vssd1 vssd1 vccd1 vccd1 _08381_ sky130_fd_sc_hd__a21boi_1
X_12979_ _05627_ _05657_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__nor2_4
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17506_ _10041_ _10042_ vssd1 vssd1 vccd1 vccd1 _10043_ sky130_fd_sc_hd__or2_1
X_14718_ _03819_ _03764_ _07333_ _05026_ rbzero.wall_tracer.wall\[1\] vssd1 vssd1
+ vccd1 vccd1 _00479_ sky130_fd_sc_hd__a32o_1
XFILLER_127_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18486_ _02231_ _02232_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__nand2_1
X_15698_ _08284_ _08311_ vssd1 vssd1 vccd1 vccd1 _08312_ sky130_fd_sc_hd__xor2_1
XFILLER_33_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17437_ _09721_ _09974_ _09852_ _09853_ vssd1 vssd1 vccd1 vccd1 _09975_ sky130_fd_sc_hd__a22o_1
XFILLER_177_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14649_ rbzero.wall_tracer.trackDistX\[6\] rbzero.wall_tracer.trackDistY\[6\] _07258_
+ vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__mux2_1
XFILLER_178_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_16 o_rgb[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_27 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_38 _10056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17368_ _09903_ _09905_ vssd1 vssd1 vccd1 vccd1 _09906_ sky130_fd_sc_hd__nand2_1
XFILLER_18_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_49 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19107_ _03808_ _02718_ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__and2_1
X_16319_ _04929_ _07652_ _08633_ vssd1 vssd1 vccd1 vccd1 _08930_ sky130_fd_sc_hd__and3_1
XFILLER_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17299_ _09706_ _09836_ _09837_ vssd1 vssd1 vccd1 vccd1 _09838_ sky130_fd_sc_hd__o21ai_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19038_ _02680_ vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21000_ net57 _01016_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_141_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20715_ net85 _00731_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20646_ net66 _00662_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20577_ net82 _00593_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_221_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10330_ rbzero.tex_r1\[59\] rbzero.tex_r1\[60\] _03366_ vssd1 vssd1 vccd1 vccd1 _03375_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10261_ rbzero.tex_b1\[28\] rbzero.tex_b1\[29\] _03333_ vssd1 vssd1 vccd1 vccd1 _03339_
+ sky130_fd_sc_hd__mux2_1
XFILLER_191_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12000_ net43 _04698_ _04708_ _04709_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__a211o_1
XFILLER_106_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10192_ rbzero.tex_b1\[61\] rbzero.tex_b1\[62\] _03300_ vssd1 vssd1 vccd1 vccd1 _03303_
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21129_ _00178_ _01145_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13951_ _06577_ _06582_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__nand2_1
XFILLER_8_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12902_ _05585_ _05590_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__nor2_2
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13882_ _06569_ _06570_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__nor2_1
X_16670_ _09254_ vssd1 vssd1 vccd1 vccd1 _09260_ sky130_fd_sc_hd__clkbuf_4
XFILLER_185_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15621_ _07377_ _07398_ _07592_ _07985_ vssd1 vssd1 vccd1 vccd1 _08235_ sky130_fd_sc_hd__or4_1
X_12833_ _05417_ _05375_ _05381_ _05372_ _05462_ _05430_ vssd1 vssd1 vccd1 vccd1 _05522_
+ sky130_fd_sc_hd__mux4_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18340_ rbzero.wall_tracer.trackDistY\[5\] rbzero.wall_tracer.stepDistY\[5\] vssd1
+ vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__and2_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _08161_ _08164_ _08165_ vssd1 vssd1 vccd1 vccd1 _08166_ sky130_fd_sc_hd__o21a_1
X_12764_ _05452_ _05428_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__xnor2_2
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ _07102_ _07184_ vssd1 vssd1 vccd1 vccd1 _07185_ sky130_fd_sc_hd__nand2_2
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11715_ rbzero.tex_g1\[40\] _04374_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__and2_1
XFILLER_203_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18271_ _02040_ _02041_ _02042_ vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__nand3_1
XFILLER_159_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15483_ _08078_ _08096_ vssd1 vssd1 vccd1 vccd1 _08097_ sky130_fd_sc_hd__xor2_1
XFILLER_30_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12695_ _05305_ _05253_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__nand2_1
XFILLER_128_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17222_ _09501_ _09503_ _09636_ _09637_ vssd1 vssd1 vccd1 vccd1 _09762_ sky130_fd_sc_hd__o31a_1
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14434_ _07105_ _07121_ vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__nand2_1
X_11646_ _04361_ _04362_ _04014_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__mux2_1
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput14 i_gpout1_sel[5] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_4
X_17153_ _09690_ _09691_ vssd1 vssd1 vccd1 vccd1 _09693_ sky130_fd_sc_hd__and2_1
Xinput25 i_gpout3_sel[4] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_4
X_14365_ _05432_ _06980_ _06984_ _06987_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__a211o_1
XFILLER_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11577_ rbzero.debug_overlay.playerX\[1\] _04234_ _04282_ rbzero.debug_overlay.playerX\[5\]
+ _04294_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__a221o_1
Xinput36 i_gpout5_sel[3] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_4
XFILLER_116_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput47 i_tex_in[0] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__buf_6
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16104_ _07519_ _08531_ vssd1 vssd1 vccd1 vccd1 _08716_ sky130_fd_sc_hd__or2_1
XFILLER_183_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13316_ _05957_ _06002_ _06003_ _06004_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__o22ai_1
X_17084_ _09446_ _09488_ _09624_ vssd1 vssd1 vccd1 vccd1 _09625_ sky130_fd_sc_hd__a21boi_1
XFILLER_183_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10528_ _03481_ vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__clkbuf_1
X_14296_ _05501_ vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__buf_2
XFILLER_170_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16035_ _08486_ _08488_ vssd1 vssd1 vccd1 vccd1 _08648_ sky130_fd_sc_hd__and2_1
X_13247_ _05879_ _05935_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__xor2_1
XFILLER_157_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10459_ _03289_ _03442_ _03443_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__or3_4
XFILLER_83_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13178_ _05859_ _05860_ _05865_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__or3_1
XFILLER_170_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12129_ net30 vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__inv_2
X_17986_ _09955_ _08663_ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__nor2_1
XFILLER_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19725_ rbzero.pov.ready_buffer\[23\] _03061_ _03063_ rbzero.debug_overlay.facingY\[-8\]
+ _03066_ vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__a221o_1
X_16937_ _09209_ _09210_ _09478_ vssd1 vssd1 vccd1 vccd1 _09479_ sky130_fd_sc_hd__a21boi_1
XFILLER_238_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19656_ _07390_ _02958_ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__nor2_1
X_16868_ _08274_ _07916_ vssd1 vssd1 vccd1 vccd1 _09410_ sky130_fd_sc_hd__nor2_1
XFILLER_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18607_ rbzero.wall_tracer.rayAddendX\[11\] _02158_ _09257_ _02344_ _02336_ vssd1
+ vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__a221o_1
X_15819_ _07788_ _08423_ _08430_ _08432_ vssd1 vssd1 vccd1 vccd1 _08433_ sky130_fd_sc_hd__o31ai_1
XFILLER_20_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19587_ rbzero.pov.ready_buffer\[62\] _07367_ _02963_ vssd1 vssd1 vccd1 vccd1 _02968_
+ sky130_fd_sc_hd__mux2_1
XFILLER_111_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16799_ rbzero.wall_tracer.trackDistX\[-4\] _09301_ _09338_ _09344_ vssd1 vssd1 vccd1
+ vccd1 _00549_ sky130_fd_sc_hd__o22a_1
XFILLER_94_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18538_ _02247_ rbzero.debug_overlay.vplaneX\[-3\] vssd1 vssd1 vccd1 vccd1 _02282_
+ sky130_fd_sc_hd__xor2_1
XFILLER_181_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18469_ rbzero.wall_tracer.rayAddendX\[0\] _00013_ _02217_ vssd1 vssd1 vccd1 vccd1
+ _00595_ sky130_fd_sc_hd__o21a_1
XFILLER_179_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20500_ net128 _00516_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20431_ net121 _00462_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20362_ _03284_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20293_ _03257_ vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__clkinv_2
XFILLER_115_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11500_ _04217_ _04207_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__and2_2
XPHY_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12480_ _05156_ _05166_ _05165_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__a21oi_1
XFILLER_138_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ rbzero.tex_r1\[39\] rbzero.tex_r1\[38\] _04148_ vssd1 vssd1 vccd1 vccd1 _04149_
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20629_ net56 _00645_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14150_ _06751_ _06779_ vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__xnor2_1
XFILLER_138_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11362_ rbzero.row_render.size\[3\] _04043_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__nand2_1
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13101_ _05616_ _05638_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__nor2_1
XFILLER_192_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10313_ _03299_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__clkbuf_4
X_14081_ _06763_ _06769_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__xor2_1
XFILLER_180_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11293_ rbzero.tex_r0\[11\] _03939_ _03941_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__and3_1
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13032_ _05688_ _05690_ _05720_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__a21o_1
XFILLER_112_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10244_ rbzero.tex_b1\[36\] rbzero.tex_b1\[37\] _03322_ vssd1 vssd1 vccd1 vccd1 _03330_
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17840_ _01619_ _01622_ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__and2_1
XFILLER_121_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10175_ gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__clkbuf_4
XTAP_6864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17771_ _01549_ _01554_ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14983_ _07519_ _07524_ vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__or2_1
XFILLER_232_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19510_ _02923_ vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16722_ _09275_ vssd1 vssd1 vccd1 vccd1 _09276_ sky130_fd_sc_hd__clkbuf_4
X_13934_ _06576_ _06622_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__xnor2_1
XFILLER_234_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19441_ rbzero.pov.spi_buffer\[18\] rbzero.pov.spi_buffer\[19\] _02877_ vssd1 vssd1
+ vccd1 vccd1 _02887_ sky130_fd_sc_hd__mux2_1
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16653_ _09252_ vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13865_ _06509_ _06536_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__xnor2_1
XFILLER_228_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15604_ _08173_ _08217_ vssd1 vssd1 vccd1 vccd1 _08218_ sky130_fd_sc_hd__nor2_1
XFILLER_62_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12816_ _05353_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__inv_2
X_19372_ _02860_ vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__clkinv_2
X_16584_ _09187_ _09192_ vssd1 vssd1 vccd1 vccd1 _09193_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13796_ _05767_ _06388_ _06422_ _06317_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__o22a_1
XFILLER_163_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18323_ _05121_ _02086_ _02087_ _02013_ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__a31o_1
XFILLER_128_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15535_ _08126_ _08128_ vssd1 vssd1 vccd1 vccd1 _08149_ sky130_fd_sc_hd__nor2_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12747_ _05391_ _05314_ _05435_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__or3_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ rbzero.wall_tracer.trackDistY\[-7\] rbzero.wall_tracer.stepDistY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__nand2_1
XFILLER_148_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15466_ _08037_ _08040_ vssd1 vssd1 vccd1 vccd1 _08080_ sky130_fd_sc_hd__xor2_1
X_12678_ _05296_ _05233_ _05263_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__and3_1
XFILLER_230_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17205_ _09619_ _09621_ vssd1 vssd1 vccd1 vccd1 _09745_ sky130_fd_sc_hd__or2b_1
XFILLER_54_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14417_ _07103_ _07104_ _07105_ vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__mux2_1
XFILLER_15_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11629_ _04344_ _04345_ _04014_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__mux2_1
X_18185_ _01846_ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__inv_2
X_15397_ _07842_ _07936_ vssd1 vssd1 vccd1 vccd1 _08011_ sky130_fd_sc_hd__nor2_1
XFILLER_184_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17136_ _09674_ _09675_ vssd1 vssd1 vccd1 vccd1 _09676_ sky130_fd_sc_hd__nor2_1
XFILLER_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14348_ _06987_ _07032_ _07033_ _07036_ _06990_ vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__o311a_1
XFILLER_171_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17067_ _07838_ _09607_ _09472_ vssd1 vssd1 vccd1 vccd1 _09608_ sky130_fd_sc_hd__and3_1
XFILLER_239_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14279_ _06688_ _06791_ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__and2_1
XFILLER_170_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16018_ _07217_ _07221_ _07225_ _07687_ _07229_ vssd1 vssd1 vccd1 vccd1 _08631_ sky130_fd_sc_hd__o41a_1
XFILLER_174_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ _01749_ _01750_ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__and2_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19708_ _03060_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__buf_2
X_20980_ net90 _00996_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19639_ _03007_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__buf_2
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20414_ net136 _00445_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21394_ net86 _01410_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20345_ _02374_ _02376_ _02375_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__a21bo_1
XFILLER_135_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20276_ _03256_ vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__clkinv_2
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ _04665_ o_rgb[7] _04689_ net19 vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__a211o_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10931_ _03692_ vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13650_ _06332_ _06334_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10862_ _03656_ vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12601_ rbzero.wall_tracer.visualWallDist\[8\] vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__clkinv_2
XFILLER_77_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13581_ _06183_ _05702_ _06269_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__and3_1
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _03620_ vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__clkbuf_1
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15320_ _07760_ _07664_ _07759_ _07761_ vssd1 vssd1 vccd1 vccd1 _07934_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_164_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12532_ _05163_ _05208_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__xnor2_4
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15251_ _07742_ _07751_ vssd1 vssd1 vccd1 vccd1 _07865_ sky130_fd_sc_hd__or2_1
XFILLER_185_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12463_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__nand2_1
XFILLER_201_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14202_ _05959_ _06423_ _06890_ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__or3b_1
XFILLER_144_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11414_ rbzero.tex_r1\[59\] _03938_ _03940_ _03915_ vssd1 vssd1 vccd1 vccd1 _04132_
+ sky130_fd_sc_hd__a31o_1
X_15182_ _07788_ _07598_ _07795_ vssd1 vssd1 vccd1 vccd1 _07796_ sky130_fd_sc_hd__or3_1
XFILLER_201_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12394_ _05044_ _05086_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__nand2_1
XFILLER_32_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14133_ _06817_ _06821_ vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11345_ rbzero.row_render.size\[6\] _03783_ _03290_ _04052_ _04063_ vssd1 vssd1 vccd1
+ vccd1 _04064_ sky130_fd_sc_hd__o221a_1
XFILLER_10_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19990_ _03121_ vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__clkinv_2
XFILLER_152_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14064_ _06740_ _06748_ _06750_ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__and3_1
XFILLER_141_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18941_ rbzero.pov.spi_buffer\[19\] rbzero.pov.ready_buffer\[19\] _02629_ vssd1 vssd1
+ vccd1 vccd1 _02630_ sky130_fd_sc_hd__mux2_1
X_11276_ rbzero.tex_r0\[27\] rbzero.tex_r0\[26\] _03936_ vssd1 vssd1 vccd1 vccd1 _03995_
+ sky130_fd_sc_hd__mux2_1
XFILLER_171_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13015_ _05566_ _05605_ _05583_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__a21o_1
X_10227_ rbzero.tex_b1\[44\] rbzero.tex_b1\[45\] _03311_ vssd1 vssd1 vccd1 vccd1 _03321_
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18872_ _02577_ _02580_ _02584_ _02586_ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__and4bb_1
XTAP_6650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17823_ _01513_ _01514_ _01606_ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__and3_1
XFILLER_132_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17754_ _10056_ _08724_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__nor2_1
XTAP_5993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14966_ _07485_ _07552_ _07553_ _07579_ vssd1 vssd1 vccd1 vccd1 _07580_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16705_ rbzero.traced_texa\[7\] _09264_ _09265_ rbzero.wall_tracer.visualWallDist\[7\]
+ vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__a22o_1
X_13917_ _06518_ _06514_ vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__nand2_1
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17685_ _01450_ _01469_ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14897_ rbzero.wall_tracer.state\[13\] rbzero.wall_tracer.stepDistY\[-10\] vssd1
+ vssd1 vccd1 vccd1 _07511_ sky130_fd_sc_hd__nand2_1
XFILLER_130_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19424_ _02878_ vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__clkbuf_1
X_16636_ _09243_ _03813_ vssd1 vssd1 vccd1 vccd1 _09244_ sky130_fd_sc_hd__nand2_2
XFILLER_78_1279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13848_ _06509_ _06536_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__and2b_1
XFILLER_63_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19355_ _02858_ vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__clkinv_2
X_16567_ _09174_ _09175_ vssd1 vssd1 vccd1 vccd1 _09176_ sky130_fd_sc_hd__xor2_1
XFILLER_16_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13779_ _06440_ _06407_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18306_ _02070_ _02071_ _02065_ _02068_ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__a211oi_1
XFILLER_31_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15518_ _08125_ _08124_ vssd1 vssd1 vccd1 vccd1 _08132_ sky130_fd_sc_hd__and2_1
XFILLER_148_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19286_ rbzero.spi_registers.new_vshift\[2\] rbzero.spi_registers.spi_buffer\[2\]
+ _02825_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__mux2_1
XFILLER_203_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16498_ rbzero.wall_tracer.texu\[4\] _07338_ _03819_ _09107_ vssd1 vssd1 vccd1 vccd1
+ _00485_ sky130_fd_sc_hd__o211a_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18237_ _01997_ _02011_ _02012_ _02013_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__a31o_1
XFILLER_198_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15449_ _07542_ _07549_ _07592_ _07985_ vssd1 vssd1 vccd1 vccd1 _08063_ sky130_fd_sc_hd__or4_1
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18168_ _09829_ _08852_ _09373_ _09833_ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__o22a_1
XFILLER_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17119_ _09652_ _09658_ vssd1 vssd1 vccd1 vccd1 _09659_ sky130_fd_sc_hd__xor2_1
XFILLER_144_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18099_ _01873_ _01878_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__or2_1
XFILLER_85_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20130_ _03093_ _03161_ _03162_ _03137_ rbzero.texV\[-7\] vssd1 vssd1 vccd1 vccd1
+ _01311_ sky130_fd_sc_hd__a32o_1
XFILLER_104_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20061_ _03129_ vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__clkinv_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20963_ net116 _00979_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20894_ net62 _00910_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21377_ _00400_ _01393_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_218_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11130_ rbzero.traced_texVinit\[3\] rbzero.spi_registers.vshift\[0\] vssd1 vssd1
+ vccd1 vccd1 _03849_ sky130_fd_sc_hd__or2_1
XFILLER_190_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20328_ gpout1.clk_div\[0\] _03003_ vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__nor2_1
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11061_ _03787_ vssd1 vssd1 vccd1 vccd1 o_tex_oeb0 sky130_fd_sc_hd__buf_4
XTAP_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20259_ _03254_ vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__clkinv_2
XTAP_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ _07429_ _07430_ _07433_ _07352_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__a22o_1
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ rbzero.debug_overlay.playerX\[-6\] _07364_ vssd1 vssd1 vccd1 vccd1 _07365_
+ sky130_fd_sc_hd__or2_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11963_ _04671_ _04672_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__or2_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _06386_ _06390_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__xnor2_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17470_ _10005_ _10007_ vssd1 vssd1 vccd1 vccd1 _10008_ sky130_fd_sc_hd__nor2_1
XFILLER_233_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10914_ rbzero.tex_b0\[41\] rbzero.tex_b0\[40\] _03682_ vssd1 vssd1 vccd1 vccd1 _03684_
+ sky130_fd_sc_hd__mux2_1
XFILLER_229_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14682_ rbzero.wall_tracer.stepDistX\[-4\] _07189_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _07315_ sky130_fd_sc_hd__mux2_1
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11894_ _03289_ _04604_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__nor2_1
XFILLER_205_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16421_ _09029_ _09030_ vssd1 vssd1 vccd1 vccd1 _09031_ sky130_fd_sc_hd__xor2_1
XFILLER_189_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13633_ _05701_ _06319_ _06321_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__and3_1
X_10845_ _03647_ vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19140_ _09243_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__clkbuf_4
XFILLER_213_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16352_ _08838_ _08962_ vssd1 vssd1 vccd1 vccd1 _08963_ sky130_fd_sc_hd__xnor2_1
X_13564_ _06250_ _06252_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__xor2_1
XFILLER_125_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10776_ _03611_ vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15303_ _07602_ _07916_ vssd1 vssd1 vccd1 vccd1 _07917_ sky130_fd_sc_hd__nor2_1
XFILLER_160_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12515_ _05200_ _05201_ _05203_ _03789_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__a22oi_4
X_19071_ rbzero.spi_registers.spi_buffer\[7\] rbzero.spi_registers.spi_buffer\[6\]
+ _02690_ vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__mux2_1
X_16283_ _07890_ _07553_ _08893_ _07726_ vssd1 vssd1 vccd1 vccd1 _08894_ sky130_fd_sc_hd__and4b_1
X_13495_ _06183_ _05850_ _05849_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__o21ba_1
XFILLER_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18022_ _09018_ _09115_ _01652_ _01653_ vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__o31a_1
XFILLER_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15234_ _07647_ _07653_ vssd1 vssd1 vccd1 vccd1 _07848_ sky130_fd_sc_hd__nand2_1
XFILLER_173_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12446_ _05136_ rbzero.map_rom.a6 _05028_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__mux2_1
XFILLER_139_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15165_ _07774_ _07778_ vssd1 vssd1 vccd1 vccd1 _07779_ sky130_fd_sc_hd__xnor2_1
X_12377_ _05067_ _05069_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__nand2_1
XFILLER_126_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14116_ _06746_ _06803_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__nand2_1
X_11328_ rbzero.row_render.size\[7\] _04046_ rbzero.row_render.size\[8\] vssd1 vssd1
+ vccd1 vccd1 _04047_ sky130_fd_sc_hd__o21a_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15096_ _07466_ rbzero.wall_tracer.stepDistX\[-1\] vssd1 vssd1 vccd1 vccd1 _07710_
+ sky130_fd_sc_hd__nand2_1
XFILLER_153_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19973_ _03120_ vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__clkinv_2
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18924_ rbzero.pov.spi_buffer\[11\] rbzero.pov.ready_buffer\[11\] _02618_ vssd1 vssd1
+ vccd1 vccd1 _02621_ sky130_fd_sc_hd__mux2_1
X_14047_ _06734_ _06735_ vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__xnor2_1
X_11259_ rbzero.tex_r0\[33\] rbzero.tex_r0\[32\] _03974_ vssd1 vssd1 vccd1 vccd1 _03978_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18855_ _02557_ _02555_ _02564_ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__and3_1
XTAP_6480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17806_ _10121_ _01589_ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__xnor2_1
XFILLER_132_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18786_ _02478_ _02487_ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__or2_1
XFILLER_227_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15998_ _08609_ _08610_ vssd1 vssd1 vccd1 vccd1 _08611_ sky130_fd_sc_hd__and2b_1
XFILLER_94_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17737_ _01445_ _01516_ _01520_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__a21o_1
X_14949_ rbzero.debug_overlay.playerX\[-2\] _07492_ rbzero.debug_overlay.playerX\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _07563_ sky130_fd_sc_hd__o21ai_1
XFILLER_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17668_ _09428_ _07827_ _09963_ _09163_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_169_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19407_ _02869_ vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_223_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16619_ _09226_ _09227_ vssd1 vssd1 vccd1 vccd1 _09228_ sky130_fd_sc_hd__xor2_1
XFILLER_211_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17599_ _10133_ _10135_ vssd1 vssd1 vccd1 vccd1 _10136_ sky130_fd_sc_hd__nor2_1
XFILLER_56_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19338_ _02855_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__buf_4
XFILLER_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19269_ rbzero.spi_registers.new_other\[6\] rbzero.spi_registers.spi_buffer\[6\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__mux2_1
XFILLER_164_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21300_ net134 _01316_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21231_ _00280_ _01247_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21162_ _00211_ _01178_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20113_ rbzero.traced_texa\[-9\] rbzero.texV\[-9\] vssd1 vssd1 vccd1 vccd1 _03148_
+ sky130_fd_sc_hd__or2_1
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21093_ _00142_ _01109_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20044_ _03127_ vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__clkinv_2
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20946_ net77 _00962_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20877_ net55 _00893_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_230_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10630_ rbzero.tex_g1\[47\] rbzero.tex_g1\[48\] _03530_ vssd1 vssd1 vccd1 vccd1 _03535_
+ sky130_fd_sc_hd__mux2_1
XFILLER_198_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10561_ _03498_ vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12300_ rbzero.wall_tracer.trackDistY\[11\] vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__inv_2
XFILLER_194_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13280_ _05955_ _05968_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__xnor2_1
XFILLER_212_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10492_ _03462_ vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12231_ _04927_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__buf_4
XFILLER_136_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12162_ _04858_ _04859_ _04868_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__a21o_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11113_ _03830_ _03831_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__nor2_1
X_16970_ _09509_ _09510_ _09363_ _09366_ vssd1 vssd1 vccd1 vccd1 _09512_ sky130_fd_sc_hd__a211oi_1
X_12093_ o_tex_oeb0 _04798_ _04799_ net47 _04800_ vssd1 vssd1 vccd1 vccd1 _04801_
+ sky130_fd_sc_hd__a221o_1
XFILLER_150_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15921_ _07792_ _07517_ _07620_ rbzero.wall_tracer.visualWallDist\[4\] vssd1 vssd1
+ vccd1 vccd1 _08535_ sky130_fd_sc_hd__or4b_1
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11044_ rbzero.othery\[2\] _03733_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__xnor2_1
XFILLER_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18640_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.wall_tracer.rayAddendY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__and2_1
XFILLER_231_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15852_ _07751_ _07736_ vssd1 vssd1 vccd1 vccd1 _08466_ sky130_fd_sc_hd__nor2_1
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14803_ _07213_ _07179_ _07346_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__a21o_1
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ _02166_ _02311_ _02312_ _02158_ rbzero.wall_tracer.rayAddendX\[7\] vssd1
+ vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__a32o_1
X_15783_ _08392_ _08396_ vssd1 vssd1 vccd1 vccd1 _08397_ sky130_fd_sc_hd__xor2_1
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12995_ _05670_ _05676_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17522_ _09921_ _10058_ vssd1 vssd1 vccd1 vccd1 _10059_ sky130_fd_sc_hd__nand2_1
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14734_ _07346_ _07347_ vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__nand2_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11946_ _04652_ _04654_ _04656_ _04653_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__a22o_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ _09735_ _09858_ _09861_ vssd1 vssd1 vccd1 vccd1 _09991_ sky130_fd_sc_hd__a21o_1
XFILLER_205_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14665_ rbzero.wall_tracer.visualWallDist\[11\] _07253_ _07306_ _07257_ vssd1 vssd1
+ vccd1 vccd1 _00453_ sky130_fd_sc_hd__o211a_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _04590_ vssd1 vssd1 vccd1 vccd1 o_rgb[23] sky130_fd_sc_hd__buf_4
XFILLER_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16404_ _08898_ _08899_ vssd1 vssd1 vccd1 vccd1 _09014_ sky130_fd_sc_hd__nor2_1
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13616_ _06304_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__buf_2
X_17384_ _09018_ _08855_ _09921_ vssd1 vssd1 vccd1 vccd1 _09922_ sky130_fd_sc_hd__a21oi_1
X_10828_ rbzero.tex_g0\[18\] rbzero.tex_g0\[17\] _03638_ vssd1 vssd1 vccd1 vccd1 _03639_
+ sky130_fd_sc_hd__mux2_1
X_14596_ rbzero.wall_tracer.trackDistX\[-10\] rbzero.wall_tracer.trackDistY\[-10\]
+ _07258_ vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__mux2_1
XFILLER_164_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19123_ rbzero.otherx\[3\] _02723_ _02731_ _02728_ vssd1 vssd1 vccd1 vccd1 _00735_
+ sky130_fd_sc_hd__o211a_1
X_16335_ _08806_ _08808_ vssd1 vssd1 vccd1 vccd1 _08946_ sky130_fd_sc_hd__nor2_1
XFILLER_201_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13547_ _06234_ _06235_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__nor2_1
XFILLER_125_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10759_ rbzero.tex_g0\[50\] rbzero.tex_g0\[49\] _03593_ vssd1 vssd1 vccd1 vccd1 _03602_
+ sky130_fd_sc_hd__mux2_1
XFILLER_173_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19054_ _02688_ vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__clkbuf_1
X_16266_ _08862_ _08876_ vssd1 vssd1 vccd1 vccd1 _08877_ sky130_fd_sc_hd__xnor2_1
XFILLER_199_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13478_ _06158_ _06160_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__xor2_1
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18005_ _01785_ _01786_ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__nand2_1
XFILLER_173_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15217_ _03795_ rbzero.wall_tracer.stepDistY\[2\] vssd1 vssd1 vccd1 vccd1 _07831_
+ sky130_fd_sc_hd__nor2_1
X_12429_ _03797_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__buf_6
X_16197_ _08806_ _08808_ vssd1 vssd1 vccd1 vccd1 _08809_ sky130_fd_sc_hd__xor2_1
XFILLER_127_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15148_ _07760_ _07664_ _07759_ _07761_ vssd1 vssd1 vccd1 vccd1 _07762_ sky130_fd_sc_hd__or4bb_1
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15079_ _07342_ _05186_ _07692_ vssd1 vssd1 vccd1 vccd1 _07693_ sky130_fd_sc_hd__a21o_1
X_19956_ _03118_ vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__clkinv_2
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18907_ rbzero.pov.spi_buffer\[3\] rbzero.pov.ready_buffer\[3\] _02608_ vssd1 vssd1
+ vccd1 vccd1 _02612_ sky130_fd_sc_hd__mux2_1
XFILLER_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19887_ _03111_ vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__clkinv_2
XFILLER_95_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18838_ rbzero.wall_tracer.rayAddendY\[8\] rbzero.wall_tracer.rayAddendY\[7\] _02509_
+ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__o21a_1
XFILLER_3_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18769_ _02479_ _02491_ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__xor2_1
XFILLER_243_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20800_ _00018_ _00816_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20731_ net103 _00747_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_212_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20662_ net67 _00678_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20593_ net97 _00609_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f2 sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21214_ _00263_ _01230_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21145_ _00194_ _01161_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21076_ _00125_ _01092_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20027_ _03126_ vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__clkinv_2
XFILLER_59_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11800_ _03954_ _04489_ _04497_ _04514_ _04026_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__a311o_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _05348_ _05356_ _05359_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__or3_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _03825_ _04444_ _04446_ _04301_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__a31o_4
XFILLER_242_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20929_ net74 _00945_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[66\] sky130_fd_sc_hd__dfxtp_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14450_ _07137_ vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__clkbuf_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11662_ _03980_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__clkbuf_4
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13401_ _06084_ _06083_ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__and2b_1
XFILLER_122_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10613_ rbzero.tex_g1\[55\] rbzero.tex_g1\[56\] _03519_ vssd1 vssd1 vccd1 vccd1 _03526_
+ sky130_fd_sc_hd__mux2_1
X_14381_ _07048_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__clkinv_2
X_11593_ rbzero.tex_g0\[27\] rbzero.tex_g0\[26\] _03935_ vssd1 vssd1 vccd1 vccd1 _04310_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16120_ _07621_ vssd1 vssd1 vccd1 vccd1 _08732_ sky130_fd_sc_hd__buf_2
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13332_ _05993_ _06019_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__nor2_1
X_10544_ _03489_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16051_ _07633_ _08662_ _08663_ vssd1 vssd1 vccd1 vccd1 _08664_ sky130_fd_sc_hd__or3_2
XFILLER_182_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13263_ _05907_ _05922_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__xor2_1
X_10475_ _03453_ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_237_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15002_ _07526_ _07528_ _07356_ vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__a21o_4
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12214_ _04889_ _04917_ _04919_ vssd1 vssd1 vccd1 vccd1 o_gpout[5] sky130_fd_sc_hd__o21a_2
X_13194_ _05820_ _05882_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__xnor2_2
XFILLER_237_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12145_ _04825_ net27 _04116_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__and3_1
X_19810_ _02863_ vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__clkinv_2
XFILLER_151_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16953_ _09159_ _09222_ _09494_ vssd1 vssd1 vccd1 vccd1 _09495_ sky130_fd_sc_hd__a21oi_1
X_12076_ _04591_ _04080_ _04628_ _04101_ net21 _04781_ vssd1 vssd1 vccd1 vccd1 _04784_
+ sky130_fd_sc_hd__mux4_1
X_19741_ rbzero.pov.ready_buffer\[13\] _03067_ _03068_ rbzero.debug_overlay.vplaneX\[-7\]
+ _03015_ vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__a221o_1
XFILLER_46_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15904_ _07424_ _07805_ _07892_ _07889_ vssd1 vssd1 vccd1 vccd1 _08518_ sky130_fd_sc_hd__o31a_1
X_11027_ rbzero.map_rom.f4 rbzero.map_rom.f3 _03751_ _03754_ vssd1 vssd1 vccd1 vccd1
+ _03755_ sky130_fd_sc_hd__a31o_1
XFILLER_237_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19672_ rbzero.debug_overlay.playerY\[0\] _07498_ vssd1 vssd1 vccd1 vccd1 _03032_
+ sky130_fd_sc_hd__or2_1
X_16884_ _09187_ _09192_ vssd1 vssd1 vccd1 vccd1 _09426_ sky130_fd_sc_hd__or2b_1
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18623_ _03798_ _02355_ _02356_ _02357_ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__a31o_1
X_15835_ _08355_ _08318_ _08445_ _08448_ vssd1 vssd1 vccd1 vccd1 _08449_ sky130_fd_sc_hd__a2bb2o_2
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18554_ _02295_ _02296_ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__xnor2_1
XFILLER_206_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15766_ _08358_ _08359_ _08374_ vssd1 vssd1 vccd1 vccd1 _08380_ sky130_fd_sc_hd__nand3_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12978_ _05661_ _05663_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__xor2_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _09927_ _09930_ _10040_ vssd1 vssd1 vccd1 vccd1 _10042_ sky130_fd_sc_hd__and3_1
XFILLER_209_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14717_ _03819_ _03756_ _07333_ _05026_ rbzero.wall_tracer.wall\[0\] vssd1 vssd1
+ vccd1 vccd1 _00478_ sky130_fd_sc_hd__a32o_1
XFILLER_75_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18485_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__or2_1
X_11929_ net14 _04639_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__nand2_1
XFILLER_233_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15697_ _08286_ _08309_ _08310_ vssd1 vssd1 vccd1 vccd1 _08311_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17436_ _09449_ _09603_ vssd1 vssd1 vccd1 vccd1 _09974_ sky130_fd_sc_hd__nor2_1
XFILLER_220_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14648_ rbzero.wall_tracer.visualWallDist\[5\] _07253_ _07293_ _07295_ _07266_ vssd1
+ vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__o221a_1
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 o_rgb[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_28 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ _09904_ vssd1 vssd1 vccd1 vccd1 _09905_ sky130_fd_sc_hd__inv_2
XFILLER_202_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_39 o_rgb[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14579_ _07244_ vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19106_ _04246_ _02717_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__nor2_1
X_16318_ _08478_ _08928_ _07835_ vssd1 vssd1 vccd1 vccd1 _08929_ sky130_fd_sc_hd__a21oi_1
XFILLER_203_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17298_ _07800_ _09451_ _09707_ vssd1 vssd1 vccd1 vccd1 _09837_ sky130_fd_sc_hd__or3_1
XFILLER_185_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19037_ rbzero.pov.spi_buffer\[65\] rbzero.pov.ready_buffer\[65\] _02673_ vssd1 vssd1
+ vccd1 vccd1 _02680_ sky130_fd_sc_hd__mux2_1
X_16249_ _07625_ _08721_ _08725_ _08719_ vssd1 vssd1 vccd1 vccd1 _08860_ sky130_fd_sc_hd__o31a_1
XFILLER_173_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19939_ _03117_ vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__clkinv_2
XFILLER_101_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20714_ net85 _00730_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20645_ net62 _00661_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20576_ net81 _00592_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ _03338_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10191_ _03302_ vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21128_ _00177_ _01144_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13950_ _06636_ _06638_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__nand2_1
X_21059_ _00108_ _01075_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12901_ _05406_ _05540_ _05588_ _05589_ _05480_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__o2111a_1
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13881_ _06567_ _06568_ _06563_ vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__o21a_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15620_ _07399_ _07985_ vssd1 vssd1 vccd1 vccd1 _08234_ sky130_fd_sc_hd__or2_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _05350_ _05353_ _05346_ _05438_ _05429_ _05501_ vssd1 vssd1 vccd1 vccd1 _05521_
+ sky130_fd_sc_hd__mux4_1
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15551_ _08115_ _08160_ vssd1 vssd1 vccd1 vccd1 _08165_ sky130_fd_sc_hd__or2_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _05359_ _05410_ _05437_ _05443_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__or4_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _07174_ _07050_ _07183_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__a21oi_4
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _02033_ _02035_ _02034_ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__o21bai_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ rbzero.tex_g1\[43\] rbzero.tex_g1\[42\] _03962_ vssd1 vssd1 vccd1 vccd1 _04430_
+ sky130_fd_sc_hd__mux2_1
XFILLER_202_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15482_ _08093_ _08094_ _08095_ vssd1 vssd1 vccd1 vccd1 _08096_ sky130_fd_sc_hd__a21oi_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12694_ _05284_ _05316_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__xnor2_2
XFILLER_124_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17221_ _09506_ _09638_ vssd1 vssd1 vccd1 vccd1 _09761_ sky130_fd_sc_hd__and2_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _06981_ _06980_ _07033_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__a21o_1
X_11645_ rbzero.tex_g0\[37\] rbzero.tex_g0\[36\] _04000_ vssd1 vssd1 vccd1 vccd1 _04362_
+ sky130_fd_sc_hd__mux2_1
XFILLER_202_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17152_ _09690_ _09691_ vssd1 vssd1 vccd1 vccd1 _09692_ sky130_fd_sc_hd__nor2_1
XFILLER_156_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14364_ _06985_ _06995_ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__or2_1
Xinput15 i_gpout2_sel[0] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_6
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11576_ rbzero.debug_overlay.playerX\[-2\] _04245_ _04243_ rbzero.debug_overlay.playerX\[0\]
+ _03821_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__a221o_1
Xinput26 i_gpout3_sel[5] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_4
Xinput37 i_gpout5_sel[4] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_4
X_16103_ _08591_ _08612_ _08714_ vssd1 vssd1 vccd1 vccd1 _08715_ sky130_fd_sc_hd__a21bo_1
Xinput48 i_tex_in[1] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_4
XFILLER_156_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13315_ _05957_ _06002_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17083_ _09485_ _09487_ vssd1 vssd1 vccd1 vccd1 _09624_ sky130_fd_sc_hd__or2b_1
XFILLER_196_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10527_ rbzero.tex_r0\[33\] rbzero.tex_r0\[32\] _03479_ vssd1 vssd1 vccd1 vccd1 _03481_
+ sky130_fd_sc_hd__mux2_1
XFILLER_196_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14295_ _06981_ _06979_ _06983_ vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__and3_1
XFILLER_155_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16034_ _08643_ _08646_ vssd1 vssd1 vccd1 vccd1 _08647_ sky130_fd_sc_hd__xor2_1
X_13246_ _05881_ _05934_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__and2_1
XFILLER_171_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10458_ _03291_ _03297_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__nand2_1
XFILLER_100_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13177_ _05859_ _05860_ _05865_ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__o21ai_1
XFILLER_112_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10389_ _03406_ vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12128_ _04591_ _04080_ _04628_ _04101_ _04820_ _04832_ vssd1 vssd1 vccd1 vccd1 _04835_
+ sky130_fd_sc_hd__mux4_1
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17985_ _07678_ _08531_ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__nor2_1
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16936_ _09389_ _09208_ vssd1 vssd1 vccd1 vccd1 _09478_ sky130_fd_sc_hd__nand2_1
X_12059_ _04717_ _04718_ o_rgb[14] _04721_ _04767_ vssd1 vssd1 vccd1 vccd1 o_gpout[0]
+ sky130_fd_sc_hd__o41a_4
X_19724_ rbzero.pov.ready_buffer\[22\] _03061_ _03063_ rbzero.debug_overlay.facingY\[-9\]
+ _03066_ vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__a221o_1
XFILLER_238_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16867_ _09407_ _09408_ vssd1 vssd1 vccd1 vccd1 _09409_ sky130_fd_sc_hd__nand2_1
XFILLER_168_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19655_ rbzero.debug_overlay.playerY\[-6\] _03016_ _03020_ _02978_ vssd1 vssd1 vccd1
+ vccd1 _00978_ sky130_fd_sc_hd__o211a_1
XFILLER_226_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15818_ _07616_ _07633_ _07847_ _08431_ vssd1 vssd1 vccd1 vccd1 _08432_ sky130_fd_sc_hd__or4_1
X_18606_ rbzero.wall_tracer.rayAddendX\[11\] _02343_ vssd1 vssd1 vccd1 vccd1 _02344_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_225_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19586_ _02956_ _02966_ _02967_ _02780_ vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__o211a_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16798_ _09279_ _09343_ _09283_ vssd1 vssd1 vccd1 vccd1 _09344_ sky130_fd_sc_hd__a21o_1
XFILLER_20_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18537_ _02279_ _02273_ _02276_ _09269_ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__a31oi_1
XFILLER_234_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15749_ _08361_ _08362_ vssd1 vssd1 vccd1 vccd1 _08363_ sky130_fd_sc_hd__and2_1
XFILLER_209_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18468_ _03819_ _02207_ _02216_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__a21o_1
XFILLER_178_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17419_ _09428_ _09955_ _08788_ _09163_ vssd1 vssd1 vccd1 vccd1 _09957_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18399_ _02146_ _02151_ _02152_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__o21ai_1
XFILLER_159_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20430_ net119 _00461_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20361_ _02727_ _03282_ _03283_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__and3_1
XFILLER_228_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20292_ _03257_ vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__clkinv_2
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11430_ _03934_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__buf_4
X_20628_ net54 _00644_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11361_ gpout0.hpos\[3\] vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__clkbuf_4
X_20559_ net130 _00575_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13100_ _05787_ _05788_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__nor2_1
X_10312_ _03365_ vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__clkbuf_1
X_14080_ _06719_ _06764_ _06765_ _06768_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__a22o_1
XFILLER_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11292_ rbzero.tex_r0\[9\] rbzero.tex_r0\[8\] _03961_ vssd1 vssd1 vccd1 vccd1 _04011_
+ sky130_fd_sc_hd__mux2_1
XFILLER_138_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13031_ _05691_ _05694_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__and2b_1
X_10243_ _03329_ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__clkbuf_1
XTAP_6810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17770_ _01552_ _01553_ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__xor2_1
XFILLER_43_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14982_ _07594_ _07595_ vssd1 vssd1 vccd1 vccd1 _07596_ sky130_fd_sc_hd__xnor2_1
XFILLER_120_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16721_ _09274_ vssd1 vssd1 vccd1 vccd1 _09275_ sky130_fd_sc_hd__clkbuf_4
XFILLER_134_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13933_ _06602_ _06620_ _06621_ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__a21boi_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19440_ _02886_ vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__clkbuf_1
X_16652_ _04206_ _09245_ _09251_ vssd1 vssd1 vccd1 vccd1 _09252_ sky130_fd_sc_hd__and3_1
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13864_ _06547_ _06552_ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15603_ _08188_ _08215_ _08216_ vssd1 vssd1 vccd1 vccd1 _08217_ sky130_fd_sc_hd__a21oi_1
X_12815_ _05501_ _05502_ _05503_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__a21oi_1
X_19371_ _02855_ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__buf_4
XFILLER_90_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16583_ _09183_ _09191_ vssd1 vssd1 vccd1 vccd1 _09192_ sky130_fd_sc_hd__xnor2_1
XFILLER_234_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13795_ _05861_ _06483_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__or2_1
XFILLER_62_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18322_ _02082_ _02083_ _02084_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__a21o_1
XFILLER_245_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15534_ _08116_ _08147_ vssd1 vssd1 vccd1 vccd1 _08148_ sky130_fd_sc_hd__xor2_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _05315_ _05317_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18253_ rbzero.wall_tracer.trackDistY\[-7\] rbzero.wall_tracer.stepDistY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__or2_1
XFILLER_124_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15465_ _08014_ _08016_ vssd1 vssd1 vccd1 vccd1 _08079_ sky130_fd_sc_hd__xnor2_2
XFILLER_163_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12677_ _05296_ _05262_ _05364_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__a21oi_2
X_17204_ _09717_ _09743_ vssd1 vssd1 vccd1 vccd1 _09744_ sky130_fd_sc_hd__xnor2_1
X_14416_ _05497_ vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__buf_2
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18184_ _01938_ _01963_ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__xnor2_1
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11628_ rbzero.tex_g0\[61\] rbzero.tex_g0\[60\] _04168_ vssd1 vssd1 vccd1 vccd1 _04345_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15396_ _08008_ _08009_ vssd1 vssd1 vccd1 vccd1 _08010_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17135_ _09672_ _09673_ vssd1 vssd1 vccd1 vccd1 _09675_ sky130_fd_sc_hd__and2_1
XFILLER_204_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14347_ _06985_ _07035_ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__or2_1
XFILLER_183_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11559_ rbzero.debug_overlay.playerY\[-5\] _04214_ _04237_ rbzero.debug_overlay.playerY\[-6\]
+ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__a22o_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17066_ _08923_ _09470_ vssd1 vssd1 vccd1 vccd1 _09607_ sky130_fd_sc_hd__nand2_1
X_14278_ _06686_ _06688_ vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16017_ _07689_ _07819_ _08475_ _07690_ vssd1 vssd1 vccd1 vccd1 _08630_ sky130_fd_sc_hd__and4_1
X_13229_ _05910_ _05916_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__xor2_1
XFILLER_143_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17968_ _01742_ _01748_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__or2_1
XFILLER_215_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19707_ rbzero.pov.ready _02721_ _02833_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__and3_1
XFILLER_22_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16919_ _08779_ _09055_ vssd1 vssd1 vccd1 vccd1 _09461_ sky130_fd_sc_hd__nand2_1
XFILLER_214_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17899_ _01668_ _01681_ vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__xnor2_1
XFILLER_168_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19638_ net40 _02954_ _02721_ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__o21ai_2
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19569_ _02953_ vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__clkbuf_1
XFILLER_230_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20413_ net130 _00444_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_181_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21393_ net108 _01409_ vssd1 vssd1 vccd1 vccd1 gpout1.clk_div\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20344_ _09257_ _02375_ _03273_ _02158_ rbzero.wall_tracer.rayAddendY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__a32o_1
XFILLER_179_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20275_ _03256_ vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__clkinv_2
XFILLER_103_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10930_ rbzero.tex_b0\[33\] rbzero.tex_b0\[32\] _03682_ vssd1 vssd1 vccd1 vccd1 _03692_
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10861_ rbzero.tex_g0\[2\] rbzero.tex_g0\[1\] _03649_ vssd1 vssd1 vccd1 vccd1 _03656_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12600_ _05281_ _05284_ _05286_ _05288_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__or4b_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _05621_ _05624_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__nand2_1
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10792_ rbzero.tex_g0\[35\] rbzero.tex_g0\[34\] _03616_ vssd1 vssd1 vccd1 vccd1 _03620_
+ sky130_fd_sc_hd__mux2_1
XFILLER_231_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12531_ _05219_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__buf_4
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15250_ _07748_ _07862_ _07863_ vssd1 vssd1 vccd1 vccd1 _07864_ sky130_fd_sc_hd__a21o_1
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12462_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__nand2_1
XFILLER_36_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14201_ _06858_ _06889_ vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__xor2_1
XFILLER_138_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11413_ rbzero.tex_r1\[58\] _03925_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__and2_1
X_15181_ _07791_ _07794_ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__nand2_1
XFILLER_172_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12393_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__nand2_1
XFILLER_201_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14132_ _06764_ _06818_ _06820_ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__a21bo_1
XFILLER_181_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11344_ rbzero.row_render.size\[6\] _03783_ _03780_ _04053_ _04062_ vssd1 vssd1 vccd1
+ vccd1 _04063_ sky130_fd_sc_hd__a221o_1
XFILLER_152_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14063_ _06709_ _06729_ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__xnor2_1
XFILLER_180_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18940_ _02607_ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__clkbuf_4
X_11275_ _03946_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__clkbuf_4
XFILLER_106_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13014_ _05591_ _05702_ _05566_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__or3b_4
XFILLER_84_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10226_ _03320_ vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18871_ rbzero.spi_registers.spi_counter\[2\] _02585_ vssd1 vssd1 vccd1 vccd1 _02586_
+ sky130_fd_sc_hd__xnor2_1
XTAP_6640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17822_ _01515_ _01605_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__xor2_1
XTAP_6673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17753_ _01534_ _01536_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__and2b_1
XTAP_5983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14965_ _07571_ _07572_ _07573_ vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__a21oi_4
XFILLER_212_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13916_ _06593_ _06598_ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__xor2_1
X_16704_ rbzero.traced_texa\[6\] _09264_ _09265_ rbzero.wall_tracer.visualWallDist\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__a22o_1
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17684_ _01451_ _01468_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__xnor2_1
X_14896_ _07466_ _07509_ vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__or2_1
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16635_ _03292_ vssd1 vssd1 vccd1 vccd1 _09243_ sky130_fd_sc_hd__clkbuf_4
XFILLER_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19423_ rbzero.pov.spi_buffer\[9\] rbzero.pov.spi_buffer\[10\] _02877_ vssd1 vssd1
+ vccd1 vccd1 _02878_ sky130_fd_sc_hd__mux2_1
X_13847_ _06521_ _06535_ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__nand2_1
XFILLER_21_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16566_ _08760_ _07712_ _09027_ _09025_ vssd1 vssd1 vccd1 vccd1 _09175_ sky130_fd_sc_hd__o31a_1
X_19354_ _02858_ vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__clkinv_2
XFILLER_91_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13778_ _06460_ _06466_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__xor2_1
XFILLER_210_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18305_ _02065_ _02068_ _02070_ _02071_ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__o211a_1
X_15517_ _08080_ _08090_ vssd1 vssd1 vccd1 vccd1 _08131_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12729_ _05367_ _05368_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__or2_1
XFILLER_31_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19285_ _02827_ vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16497_ _09105_ _09106_ _04933_ vssd1 vssd1 vccd1 vccd1 _09107_ sky130_fd_sc_hd__a21o_1
XFILLER_148_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18236_ _02000_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__clkbuf_4
X_15448_ _07549_ _07986_ vssd1 vssd1 vccd1 vccd1 _08062_ sky130_fd_sc_hd__or2_1
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18167_ _01768_ _01862_ _01946_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a21oi_1
XFILLER_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15379_ _07509_ _07633_ _07991_ vssd1 vssd1 vccd1 vccd1 _07993_ sky130_fd_sc_hd__o21ai_1
XFILLER_89_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17118_ _09656_ _09657_ vssd1 vssd1 vccd1 vccd1 _09658_ sky130_fd_sc_hd__nand2_1
XFILLER_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18098_ _01873_ _01878_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__nand2_1
XFILLER_172_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17049_ _09182_ _08780_ _09454_ _09452_ vssd1 vssd1 vccd1 vccd1 _09590_ sky130_fd_sc_hd__o31ai_1
XFILLER_172_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20060_ _03129_ vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__clkinv_2
XFILLER_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20962_ net91 _00978_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20893_ net62 _00909_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_246_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21376_ _00399_ _01392_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20327_ _03263_ vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11060_ _03781_ _03782_ _03785_ _03786_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__a211o_1
XFILLER_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20258_ _03254_ vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__clkinv_2
XFILLER_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20189_ rbzero.traced_texa\[3\] rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1 _03212_
+ sky130_fd_sc_hd__nand2_1
XFILLER_131_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ rbzero.debug_overlay.playerX\[-7\] rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__or3_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11962_ _04078_ _03781_ _03784_ _03291_ _04665_ _04664_ vssd1 vssd1 vccd1 vccd1 _04672_
+ sky130_fd_sc_hd__mux4_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13701_ _06317_ _06343_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__nor2_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10913_ _03683_ vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14681_ _07314_ vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__clkbuf_1
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ _04603_ _04604_ _04605_ _04080_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a31o_1
XFILLER_229_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16420_ _08896_ _08897_ _08894_ vssd1 vssd1 vccd1 vccd1 _09030_ sky130_fd_sc_hd__a21oi_1
X_13632_ _06320_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__buf_2
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10844_ rbzero.tex_g0\[10\] rbzero.tex_g0\[9\] _03638_ vssd1 vssd1 vccd1 vccd1 _03647_
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16351_ _08959_ _08961_ vssd1 vssd1 vccd1 vccd1 _08962_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13563_ _06195_ _06206_ _06251_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__a21oi_1
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10775_ rbzero.tex_g0\[43\] rbzero.tex_g0\[42\] _03605_ vssd1 vssd1 vccd1 vccd1 _03611_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15302_ _07915_ vssd1 vssd1 vccd1 vccd1 _07916_ sky130_fd_sc_hd__buf_2
XFILLER_73_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12514_ _05180_ _05202_ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__xnor2_4
X_19070_ _02697_ vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__clkbuf_1
X_16282_ _07672_ _07673_ vssd1 vssd1 vccd1 vccd1 _08893_ sky130_fd_sc_hd__nand2_1
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13494_ _05847_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__inv_2
XFILLER_125_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18021_ _01683_ _01649_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__or2b_1
XFILLER_139_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15233_ _07664_ vssd1 vssd1 vccd1 vccd1 _07847_ sky130_fd_sc_hd__clkbuf_4
XFILLER_201_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12445_ rbzero.debug_overlay.playerY\[3\] _05135_ _03798_ vssd1 vssd1 vccd1 vccd1
+ _05136_ sky130_fd_sc_hd__mux2_1
XFILLER_185_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15164_ _07775_ _07777_ vssd1 vssd1 vccd1 vccd1 _07778_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12376_ _05068_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__buf_2
XFILLER_181_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14115_ _06313_ _06634_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__nor2_1
XFILLER_126_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11327_ rbzero.row_render.size\[6\] _04045_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__and2_1
XFILLER_113_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15095_ _07708_ vssd1 vssd1 vccd1 vccd1 _07709_ sky130_fd_sc_hd__clkbuf_4
X_19972_ _03120_ vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__clkinv_2
XFILLER_119_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14046_ _05740_ _06389_ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__nor2_1
XFILLER_171_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18923_ _02620_ vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11258_ _03975_ _03976_ _03930_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__mux2_1
XFILLER_84_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10209_ rbzero.tex_b1\[53\] rbzero.tex_b1\[54\] _03311_ vssd1 vssd1 vccd1 vccd1 _03312_
+ sky130_fd_sc_hd__mux2_1
XFILLER_228_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18854_ rbzero.wall_tracer.rayAddendY\[10\] rbzero.wall_tracer.rayAddendY\[9\] _02556_
+ _02510_ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__or4b_1
XFILLER_228_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11189_ _03860_ _03894_ _03907_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__nor3b_4
XTAP_6481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17805_ _01584_ _01588_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__xor2_1
XFILLER_227_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15997_ _08607_ _08608_ vssd1 vssd1 vccd1 vccd1 _08610_ sky130_fd_sc_hd__nand2_1
XFILLER_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18785_ _02505_ _02506_ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__nand2_1
XTAP_5780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17736_ _01518_ _01519_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__nand2_1
X_14948_ rbzero.debug_overlay.playerX\[-1\] rbzero.debug_overlay.playerX\[-2\] _07492_
+ vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__or3_1
XFILLER_76_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17667_ _08067_ _09428_ _07827_ _09451_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__or4_1
X_14879_ rbzero.debug_overlay.playerX\[-2\] vssd1 vssd1 vccd1 vccd1 _07493_ sky130_fd_sc_hd__inv_2
XFILLER_51_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19406_ rbzero.pov.spi_buffer\[1\] rbzero.pov.spi_buffer\[2\] _02866_ vssd1 vssd1
+ vccd1 vccd1 _02869_ sky130_fd_sc_hd__mux2_1
X_16618_ _08974_ _09088_ _09087_ vssd1 vssd1 vccd1 vccd1 _09227_ sky130_fd_sc_hd__a21boi_1
XFILLER_63_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17598_ _09950_ _10004_ _10134_ vssd1 vssd1 vccd1 vccd1 _10135_ sky130_fd_sc_hd__a21oi_1
XFILLER_211_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16549_ _09156_ _09157_ vssd1 vssd1 vccd1 vccd1 _09158_ sky130_fd_sc_hd__nand2_1
XFILLER_204_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19337_ _02856_ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__clkinv_2
XFILLER_204_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19268_ _02818_ vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18219_ rbzero.wall_tracer.trackDistY\[-12\] rbzero.wall_tracer.stepDistY\[-12\]
+ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__nand2_1
XFILLER_163_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19199_ rbzero.spi_registers.new_vshift\[3\] _02775_ vssd1 vssd1 vccd1 vccd1 _02779_
+ sky130_fd_sc_hd__or2_1
XFILLER_129_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21230_ _00279_ _01246_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21161_ _00210_ _01177_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20112_ rbzero.texV\[-10\] _02989_ _03142_ _03147_ vssd1 vssd1 vccd1 vccd1 _01308_
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21092_ _00141_ _01108_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20043_ _03127_ vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__clkinv_2
XFILLER_115_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20945_ net77 _00961_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20876_ net58 _00892_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10560_ rbzero.tex_r0\[17\] rbzero.tex_r0\[16\] _03490_ vssd1 vssd1 vccd1 vccd1 _03498_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10491_ rbzero.tex_r0\[50\] rbzero.tex_r0\[49\] _03457_ vssd1 vssd1 vccd1 vccd1 _03462_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12230_ rbzero.wall_tracer.state\[6\] vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__inv_2
XFILLER_136_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12161_ _04836_ net29 _04864_ _04867_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__a31o_1
XFILLER_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21359_ _00382_ _01375_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11112_ rbzero.traced_texVinit\[7\] rbzero.spi_registers.vshift\[4\] vssd1 vssd1
+ vccd1 vccd1 _03831_ sky130_fd_sc_hd__nor2_1
XFILLER_151_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12092_ net48 _04773_ _04768_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__and3_1
XFILLER_81_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15920_ _08533_ vssd1 vssd1 vccd1 vccd1 _08534_ sky130_fd_sc_hd__inv_2
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11043_ rbzero.othery\[3\] _03744_ rbzero.map_rom.i_row\[4\] _03766_ _03770_ vssd1
+ vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__a221o_1
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15851_ _07862_ _08463_ _08464_ vssd1 vssd1 vccd1 vccd1 _08465_ sky130_fd_sc_hd__o21ai_1
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _04936_ _07409_ _07415_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__o21ai_4
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15782_ _07788_ _07843_ _08394_ _08395_ vssd1 vssd1 vccd1 vccd1 _08396_ sky130_fd_sc_hd__o31a_1
X_18570_ _02309_ _02310_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__or2_1
XFILLER_224_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12994_ _05678_ _05680_ _05681_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__a21o_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17521_ _10056_ _08985_ vssd1 vssd1 vccd1 vccd1 _10058_ sky130_fd_sc_hd__nor2_1
X_14733_ _05085_ _05226_ _07341_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__mux2_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11945_ net51 _04643_ _04644_ net53 _04655_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__a221o_1
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _09733_ _09735_ _09988_ vssd1 vssd1 vccd1 vccd1 _09990_ sky130_fd_sc_hd__nand3_1
XFILLER_206_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14664_ rbzero.wall_tracer.trackDistY\[11\] rbzero.wall_tracer.trackDistX\[11\] _03799_
+ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__a21o_1
XFILLER_45_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11876_ _03826_ _04589_ _04301_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__o21ba_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ _08975_ _09012_ vssd1 vssd1 vccd1 vccd1 _09013_ sky130_fd_sc_hd__xnor2_1
XFILLER_220_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13615_ _06260_ _06289_ _06303_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17383_ rbzero.wall_tracer.visualWallDist\[6\] _03796_ _08123_ vssd1 vssd1 vccd1
+ vccd1 _09921_ sky130_fd_sc_hd__and3_1
XFILLER_158_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10827_ _03604_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__clkbuf_4
X_14595_ _05025_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__buf_4
XFILLER_220_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16334_ _08903_ _08944_ vssd1 vssd1 vccd1 vccd1 _08945_ sky130_fd_sc_hd__xor2_1
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19122_ rbzero.spi_registers.new_other\[9\] _02725_ vssd1 vssd1 vccd1 vccd1 _02731_
+ sky130_fd_sc_hd__or2_1
XFILLER_186_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13546_ _06186_ _06187_ _06233_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__nor3_1
XFILLER_203_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10758_ _03601_ vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19053_ rbzero.pov.spi_buffer\[73\] rbzero.pov.ready_buffer\[73\] _02607_ vssd1 vssd1
+ vccd1 vccd1 _02688_ sky130_fd_sc_hd__mux2_1
X_16265_ _08874_ _08875_ vssd1 vssd1 vccd1 vccd1 _08876_ sky130_fd_sc_hd__nor2_1
XFILLER_145_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13477_ _06161_ _06163_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__xor2_1
X_10689_ rbzero.tex_g1\[19\] rbzero.tex_g1\[20\] _03563_ vssd1 vssd1 vccd1 vccd1 _03566_
+ sky130_fd_sc_hd__mux2_1
X_18004_ _10095_ _08735_ _01784_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__o21ai_1
X_15216_ _07815_ _07829_ vssd1 vssd1 vccd1 vccd1 _07830_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12428_ _05120_ vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16196_ _08626_ _08652_ _08807_ vssd1 vssd1 vccd1 vccd1 _08808_ sky130_fd_sc_hd__a21oi_1
X_15147_ _07675_ _07709_ _07735_ _07646_ vssd1 vssd1 vccd1 vccd1 _07761_ sky130_fd_sc_hd__o22ai_1
X_12359_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] _05050_
+ _05051_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__a211o_1
XFILLER_114_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15078_ _07334_ _05069_ _05112_ _04932_ vssd1 vssd1 vccd1 vccd1 _07692_ sky130_fd_sc_hd__a31o_1
X_19955_ _03118_ vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__clkinv_2
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14029_ _06670_ _06668_ _06516_ vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__a21o_1
X_18906_ _02611_ vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__clkbuf_1
X_19886_ _03111_ vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__clkinv_2
XFILLER_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18837_ _02533_ _02544_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__and2b_1
XFILLER_83_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18768_ _02428_ rbzero.debug_overlay.vplaneY\[-4\] vssd1 vssd1 vccd1 vccd1 _02491_
+ sky130_fd_sc_hd__xor2_1
XFILLER_208_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17719_ _01500_ _01503_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__or2_1
XFILLER_222_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18699_ _02287_ _02420_ _02421_ _02426_ vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__a31o_1
XFILLER_63_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20730_ net100 _00746_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20661_ net67 _00677_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20592_ net97 _00608_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f3 sky130_fd_sc_hd__dfxtp_2
XFILLER_108_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21213_ _00262_ _01229_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21144_ _00193_ _01160_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21075_ _00124_ _01091_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20026_ _03125_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__buf_4
XFILLER_150_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _04099_ _04445_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__nand2_1
XFILLER_226_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20928_ net75 _00944_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[65\] sky130_fd_sc_hd__dfxtp_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11661_ _04375_ _04376_ _03968_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__mux2_1
XFILLER_230_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20859_ _00077_ _00875_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13400_ _06068_ _06088_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__or2b_1
X_10612_ _03525_ vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__clkbuf_1
X_14380_ _07029_ _07064_ _07065_ _07068_ vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__a31o_1
XFILLER_161_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11592_ _04305_ _04308_ _03923_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__mux2_1
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13331_ _05993_ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__xor2_1
XFILLER_35_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10543_ rbzero.tex_r0\[25\] rbzero.tex_r0\[24\] _03479_ vssd1 vssd1 vccd1 vccd1 _03489_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16050_ rbzero.wall_tracer.visualWallDist\[7\] _03796_ vssd1 vssd1 vccd1 vccd1 _08663_
+ sky130_fd_sc_hd__nand2_2
XFILLER_155_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13262_ _05947_ _05938_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__xnor2_1
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10474_ rbzero.tex_r0\[58\] rbzero.tex_r0\[57\] _03446_ vssd1 vssd1 vccd1 vccd1 _03453_
+ sky130_fd_sc_hd__mux2_1
X_15001_ _07590_ _07614_ vssd1 vssd1 vccd1 vccd1 _07615_ sky130_fd_sc_hd__or2b_1
XFILLER_237_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12213_ _04918_ o_rgb[23] _04885_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__or3b_1
XFILLER_68_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13193_ _05705_ _05819_ _05821_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__o21bai_1
XFILLER_194_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12144_ o_tex_oeb0 _04848_ _04849_ net47 _04850_ vssd1 vssd1 vccd1 vccd1 _04851_
+ sky130_fd_sc_hd__a221o_1
XFILLER_155_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19740_ rbzero.pov.ready_buffer\[12\] _03067_ _03068_ rbzero.debug_overlay.vplaneX\[-8\]
+ _03066_ vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__a221o_1
X_16952_ _09220_ _09221_ vssd1 vssd1 vccd1 vccd1 _09494_ sky130_fd_sc_hd__nor2_1
X_12075_ _04781_ _04782_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__or2_1
XFILLER_238_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15903_ _08515_ _08516_ vssd1 vssd1 vccd1 vccd1 _08517_ sky130_fd_sc_hd__xnor2_1
X_11026_ rbzero.map_rom.f4 rbzero.map_rom.d6 _03740_ _03753_ vssd1 vssd1 vccd1 vccd1
+ _03754_ sky130_fd_sc_hd__o31ai_1
X_19671_ rbzero.debug_overlay.playerY\[-1\] _03016_ _03030_ _03031_ vssd1 vssd1 vccd1
+ vccd1 _00983_ sky130_fd_sc_hd__o211a_1
XFILLER_81_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16883_ _09168_ _09176_ _09424_ vssd1 vssd1 vccd1 vccd1 _09425_ sky130_fd_sc_hd__a21o_1
XFILLER_237_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18622_ rbzero.debug_overlay.playerX\[2\] _04940_ vssd1 vssd1 vccd1 vccd1 _02357_
+ sky130_fd_sc_hd__and2_1
XFILLER_65_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15834_ _08318_ _08447_ vssd1 vssd1 vccd1 vccd1 _08448_ sky130_fd_sc_hd__xnor2_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18553_ _02261_ _02282_ _02285_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a21o_1
X_15765_ _08377_ _08378_ vssd1 vssd1 vccd1 vccd1 _08379_ sky130_fd_sc_hd__nor2_1
X_12977_ _05650_ _05665_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__xnor2_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17504_ _09927_ _09930_ _10040_ vssd1 vssd1 vccd1 vccd1 _10041_ sky130_fd_sc_hd__a21oi_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14716_ _07332_ _03777_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__nor2_1
X_11928_ _04630_ net11 vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__nor2_1
XFILLER_244_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15696_ _08287_ _08308_ vssd1 vssd1 vccd1 vccd1 _08310_ sky130_fd_sc_hd__nor2_1
X_18484_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__nand2_1
XFILLER_178_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17435_ _09952_ _09972_ vssd1 vssd1 vccd1 vccd1 _09973_ sky130_fd_sc_hd__xor2_1
X_14647_ _07294_ _07246_ _07249_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__o21ai_1
XFILLER_177_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11859_ rbzero.tex_b1\[9\] rbzero.tex_b1\[8\] _04544_ vssd1 vssd1 vccd1 vccd1 _04573_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_18 o_rgb[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17366_ _07882_ _09115_ _09792_ _09793_ vssd1 vssd1 vccd1 vccd1 _09904_ sky130_fd_sc_hd__o31a_1
X_14578_ rbzero.wall_tracer.stepDistY\[11\] _07243_ _04925_ vssd1 vssd1 vccd1 vccd1
+ _07244_ sky130_fd_sc_hd__mux2_1
XANTENNA_29 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19105_ _02716_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__inv_2
XFILLER_14_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16317_ _04937_ rbzero.wall_tracer.stepDistX\[6\] vssd1 vssd1 vccd1 vccd1 _08928_
+ sky130_fd_sc_hd__nand2_2
X_13529_ _06177_ _06217_ vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17297_ _08240_ _09451_ vssd1 vssd1 vccd1 vccd1 _09836_ sky130_fd_sc_hd__nor2_1
XFILLER_186_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16248_ _08857_ _08858_ vssd1 vssd1 vccd1 vccd1 _08859_ sky130_fd_sc_hd__xnor2_1
X_19036_ _02679_ vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16179_ _08779_ _08636_ _08786_ _08789_ vssd1 vssd1 vccd1 vccd1 _08791_ sky130_fd_sc_hd__a22o_1
XFILLER_127_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19938_ _03117_ vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__clkinv_2
XFILLER_25_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19869_ _03109_ vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__clkinv_2
XFILLER_25_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20713_ net109 _00729_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20644_ net66 _00660_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20575_ net81 _00591_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_221_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10190_ rbzero.tex_b1\[62\] rbzero.tex_b1\[63\] _03300_ vssd1 vssd1 vccd1 vccd1 _03302_
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21127_ _00176_ _01143_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21058_ _00107_ _01074_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_219_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12900_ _05253_ _05458_ _05501_ _05431_ _05407_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__a41o_1
XFILLER_19_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20009_ _03123_ vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__clkinv_2
XFILLER_246_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13880_ _06563_ _06567_ _06568_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__nor3_1
XFILLER_41_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12831_ _05499_ _05519_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__or2_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15550_ _08162_ _08157_ _08163_ vssd1 vssd1 vccd1 vccd1 _08164_ sky130_fd_sc_hd__a21oi_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _05450_ _05343_ _05448_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__mux2_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14501_ _07107_ _07149_ _07182_ vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__a21oi_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11713_ _03958_ _04426_ _04427_ _04428_ _03924_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__o221a_1
XFILLER_163_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15481_ _08079_ _08092_ vssd1 vssd1 vccd1 vccd1 _08095_ sky130_fd_sc_hd__and2b_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _05376_ _05379_ _05381_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__or3_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _09757_ _09759_ vssd1 vssd1 vccd1 vccd1 _09760_ sky130_fd_sc_hd__nand2_2
XFILLER_187_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14432_ _05432_ _06993_ _07032_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__a21oi_1
XFILLER_159_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11644_ rbzero.tex_g0\[39\] rbzero.tex_g0\[38\] _04000_ vssd1 vssd1 vccd1 vccd1 _04361_
+ sky130_fd_sc_hd__mux2_1
XFILLER_230_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17151_ _09546_ _09555_ _09553_ vssd1 vssd1 vccd1 vccd1 _09691_ sky130_fd_sc_hd__a21oi_1
XFILLER_196_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14363_ _07007_ _07038_ _07051_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__o21ai_1
XFILLER_195_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput16 i_gpout2_sel[1] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_8
X_11575_ rbzero.debug_overlay.playerX\[-8\] _04218_ _04238_ rbzero.debug_overlay.playerX\[-7\]
+ _04292_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__a221o_1
XFILLER_122_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput27 i_gpout4_sel[0] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_6
XFILLER_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16102_ _08613_ _08590_ vssd1 vssd1 vccd1 vccd1 _08714_ sky130_fd_sc_hd__or2b_1
XFILLER_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13314_ _05607_ _05660_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__or2_1
Xinput38 i_gpout5_sel[5] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_6
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17082_ _09589_ _09622_ vssd1 vssd1 vccd1 vccd1 _09623_ sky130_fd_sc_hd__xnor2_1
X_10526_ _03480_ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__clkbuf_1
Xinput49 i_tex_in[2] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_4
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14294_ _06402_ _06982_ _06976_ _06371_ vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__o211ai_1
XFILLER_171_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16033_ _07843_ _08645_ vssd1 vssd1 vccd1 vccd1 _08646_ sky130_fd_sc_hd__nor2_1
XFILLER_171_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13245_ _05932_ _05933_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__and2b_1
XFILLER_196_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10457_ net46 net45 vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__xnor2_4
XFILLER_237_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13176_ _05862_ _05864_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__xnor2_1
X_10388_ rbzero.tex_r1\[32\] rbzero.tex_r1\[33\] _03400_ vssd1 vssd1 vccd1 vccd1 _03406_
+ sky130_fd_sc_hd__mux2_1
XFILLER_233_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12127_ _04832_ _04833_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__or2_1
XFILLER_112_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17984_ _01764_ _01765_ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__xnor2_1
X_19723_ rbzero.pov.ready_buffer\[43\] _03061_ _03063_ rbzero.debug_overlay.facingX\[10\]
+ _03066_ vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__a221o_1
X_16935_ _09201_ _09473_ _09476_ vssd1 vssd1 vccd1 vccd1 _09477_ sky130_fd_sc_hd__o21ba_1
XFILLER_238_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12058_ _04729_ _04746_ _04752_ _04766_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__or4_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11009_ _03736_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__inv_2
XFILLER_38_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19654_ rbzero.pov.ready_buffer\[47\] _02836_ _03008_ _03019_ vssd1 vssd1 vccd1 vccd1
+ _03020_ sky130_fd_sc_hd__a211o_1
X_16866_ _08086_ _07621_ _08536_ _08135_ vssd1 vssd1 vccd1 vccd1 _09408_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18605_ _02341_ _02275_ _02342_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__mux2_1
XFILLER_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15817_ _07788_ _07680_ _08389_ vssd1 vssd1 vccd1 vccd1 _08431_ sky130_fd_sc_hd__a21oi_1
X_19585_ _07462_ _02960_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__nand2_1
XFILLER_80_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16797_ _09341_ _09342_ vssd1 vssd1 vccd1 vccd1 _09343_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18536_ _02273_ _02276_ _02279_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__a21o_1
X_15748_ _08296_ _07971_ _07986_ _07470_ vssd1 vssd1 vccd1 vccd1 _08362_ sky130_fd_sc_hd__o22ai_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18467_ _03729_ _02214_ _02215_ _02197_ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__a31o_1
X_15679_ _07466_ _07675_ vssd1 vssd1 vccd1 vccd1 _08293_ sky130_fd_sc_hd__nor2_1
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17418_ _08594_ _09428_ _09955_ _08780_ vssd1 vssd1 vccd1 vccd1 _09956_ sky130_fd_sc_hd__or4_1
XFILLER_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18398_ rbzero.debug_overlay.vplaneX\[-7\] rbzero.wall_tracer.rayAddendX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__nand2_1
XFILLER_18_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17349_ _09345_ _09887_ vssd1 vssd1 vccd1 vccd1 _09888_ sky130_fd_sc_hd__and2_1
XFILLER_53_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20360_ gpout3.clk_div\[1\] gpout3.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__or2_1
XFILLER_105_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19019_ _02670_ vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20291_ _03257_ vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__clkinv_2
XFILLER_179_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20627_ net54 _00643_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11360_ rbzero.row_render.size\[4\] _04044_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20558_ net136 _00574_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10311_ rbzero.tex_b1\[4\] rbzero.tex_b1\[5\] _03355_ vssd1 vssd1 vccd1 vccd1 _03365_
+ sky130_fd_sc_hd__mux2_1
X_11291_ _04008_ _04009_ _03930_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__mux2_1
XFILLER_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20489_ net112 _00505_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_238_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13030_ _05712_ _05718_ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__nand2_1
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10242_ rbzero.tex_b1\[37\] rbzero.tex_b1\[38\] _03322_ vssd1 vssd1 vccd1 vccd1 _03329_
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14981_ _07509_ _07529_ vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__nor2_1
XTAP_6899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16720_ _09273_ vssd1 vssd1 vccd1 vccd1 _09274_ sky130_fd_sc_hd__buf_4
XFILLER_134_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13932_ _06619_ _06604_ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__or2b_1
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13863_ _06548_ _06551_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__xnor2_1
X_16651_ _03294_ _04205_ vssd1 vssd1 vccd1 vccd1 _09251_ sky130_fd_sc_hd__or2_1
XFILLER_78_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12814_ _05253_ _05462_ _05463_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__and3_1
X_15602_ _08189_ _08214_ vssd1 vssd1 vccd1 vccd1 _08216_ sky130_fd_sc_hd__nor2_1
XFILLER_90_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19370_ _02859_ vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__clkinv_2
X_16582_ _09047_ _09188_ _09189_ _09190_ vssd1 vssd1 vccd1 vccd1 _09191_ sky130_fd_sc_hd__o22a_1
X_13794_ _06482_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__buf_2
XFILLER_234_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18321_ _02085_ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__inv_2
XFILLER_231_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12745_ _05433_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__buf_4
X_15533_ _08130_ _08145_ _08146_ vssd1 vssd1 vccd1 vccd1 _08147_ sky130_fd_sc_hd__a21oi_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15464_ _08076_ _08077_ vssd1 vssd1 vccd1 vccd1 _08078_ sky130_fd_sc_hd__or2_1
X_18252_ rbzero.wall_tracer.trackDistY\[-8\] _01996_ _02026_ _09310_ vssd1 vssd1 vccd1
+ vccd1 _00569_ sky130_fd_sc_hd__o22a_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12676_ _05295_ _05364_ _05262_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__and3_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17203_ _09740_ _09742_ vssd1 vssd1 vccd1 vccd1 _09743_ sky130_fd_sc_hd__xnor2_1
X_14415_ _05432_ _06992_ _06984_ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__a21o_1
XFILLER_175_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11627_ rbzero.tex_g0\[63\] rbzero.tex_g0\[62\] _04168_ vssd1 vssd1 vccd1 vccd1 _04344_
+ sky130_fd_sc_hd__mux2_1
X_18183_ _01939_ _01962_ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__xnor2_1
X_15395_ _07439_ _07440_ _07718_ vssd1 vssd1 vccd1 vccd1 _08009_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17134_ _09672_ _09673_ vssd1 vssd1 vccd1 vccd1 _09674_ sky130_fd_sc_hd__nor2_1
XFILLER_204_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14346_ _05432_ _06993_ _07034_ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__a21o_1
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11558_ _04104_ _04106_ _04251_ _04275_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17065_ _09604_ _09605_ vssd1 vssd1 vccd1 vccd1 _09606_ sky130_fd_sc_hd__and2_1
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10509_ _03471_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__clkbuf_1
X_14277_ _06788_ _06841_ _06962_ _06964_ _06965_ vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__a221o_1
XFILLER_195_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11489_ _03293_ _04204_ _04206_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__o21ai_4
XFILLER_48_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16016_ _07453_ vssd1 vssd1 vccd1 vccd1 _08629_ sky130_fd_sc_hd__clkbuf_4
XFILLER_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13228_ _05910_ _05916_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__and2b_1
XFILLER_131_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13159_ _05624_ _05749_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__nor2_1
XFILLER_135_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _01742_ _01748_ vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__nand2_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19706_ rbzero.pov.ready_buffer\[33\] _03056_ _03059_ rbzero.debug_overlay.facingX\[-9\]
+ _03031_ vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__o221a_1
X_16918_ _09448_ _09459_ vssd1 vssd1 vccd1 vccd1 _09460_ sky130_fd_sc_hd__xor2_1
XFILLER_226_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17898_ _01678_ _01680_ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__xor2_1
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19637_ _03004_ _03006_ _03003_ vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__a21o_1
XFILLER_93_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16849_ _09387_ _09390_ vssd1 vssd1 vccd1 vccd1 _09391_ sky130_fd_sc_hd__xor2_1
XFILLER_81_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19568_ rbzero.pov.sclk_buffer\[2\] rbzero.pov.sclk_buffer\[1\] _09243_ vssd1 vssd1
+ vccd1 vccd1 _02953_ sky130_fd_sc_hd__mux2_1
XFILLER_168_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18519_ _02191_ rbzero.debug_overlay.vplaneX\[-5\] _02261_ _02262_ vssd1 vssd1 vccd1
+ vccd1 _02264_ sky130_fd_sc_hd__or4_1
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19499_ _02917_ vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20412_ net130 _00443_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_105_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21392_ net114 _01408_ vssd1 vssd1 vccd1 vccd1 gpout1.clk_div\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20343_ rbzero.debug_overlay.vplaneY\[-9\] rbzero.wall_tracer.rayAddendY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__or2_1
XFILLER_107_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20274_ _03256_ vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__clkinv_2
XTAP_6107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10860_ _03655_ vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10791_ _03619_ vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__clkbuf_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12530_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__inv_2
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12461_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__nor2_1
XFILLER_138_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14200_ _06101_ _06541_ vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__or2_1
X_11412_ rbzero.tex_r1\[57\] rbzero.tex_r1\[56\] _03935_ vssd1 vssd1 vccd1 vccd1 _04130_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15180_ _07792_ _07790_ _07579_ _07793_ vssd1 vssd1 vccd1 vccd1 _07794_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_197_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12392_ _05036_ _05082_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__xor2_2
XFILLER_240_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14131_ _05959_ _06343_ _06819_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__or3b_1
X_11343_ _04053_ _03780_ gpout0.hpos\[4\] _04054_ _04061_ vssd1 vssd1 vccd1 vccd1
+ _04062_ sky130_fd_sc_hd__o221a_1
XFILLER_193_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14062_ _06740_ _06748_ _06750_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__a21oi_2
XFILLER_158_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11274_ _03989_ _03992_ _03924_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__mux2_1
XFILLER_98_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13013_ _05604_ _05582_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__or2_1
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10225_ rbzero.tex_b1\[45\] rbzero.tex_b1\[46\] _03311_ vssd1 vssd1 vccd1 vccd1 _03320_
+ sky130_fd_sc_hd__mux2_1
XFILLER_133_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18870_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[0\] _02579_
+ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__a21o_1
XTAP_6630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17821_ _01603_ _01604_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__xnor2_1
XFILLER_132_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17752_ _09571_ _08717_ _01535_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__or3_1
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14964_ _07485_ _07542_ _07550_ _07575_ vssd1 vssd1 vccd1 vccd1 _07578_ sky130_fd_sc_hd__or4_1
XTAP_5984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16703_ rbzero.traced_texa\[5\] _09264_ _09265_ rbzero.wall_tracer.visualWallDist\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__a22o_1
X_13915_ _06535_ _06603_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__and2_1
XFILLER_48_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17683_ _01457_ _01467_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__xor2_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14895_ rbzero.wall_tracer.visualWallDist\[1\] _03795_ vssd1 vssd1 vccd1 vccd1 _07509_
+ sky130_fd_sc_hd__nand2_4
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19422_ _02865_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__clkbuf_4
XFILLER_207_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16634_ _04933_ _09241_ _09242_ _07257_ vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__o211a_1
X_13846_ _06532_ _06533_ _06534_ vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__or3_1
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19353_ _02858_ vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__clkinv_2
X_16565_ _09169_ _09173_ vssd1 vssd1 vccd1 vccd1 _09174_ sky130_fd_sc_hd__xnor2_1
X_13777_ _06462_ _06465_ vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__and2_1
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10989_ rbzero.tex_b0\[5\] rbzero.tex_b0\[4\] _03715_ vssd1 vssd1 vccd1 vccd1 _03723_
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18304_ rbzero.wall_tracer.trackDistY\[0\] rbzero.wall_tracer.stepDistY\[0\] vssd1
+ vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__nand2_1
XFILLER_71_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15516_ _08121_ _08129_ vssd1 vssd1 vccd1 vccd1 _08130_ sky130_fd_sc_hd__xor2_1
XFILLER_188_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12728_ _05365_ _05366_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__nor2_4
XFILLER_128_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19284_ rbzero.spi_registers.new_vshift\[1\] rbzero.spi_registers.spi_buffer\[1\]
+ _02825_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__mux2_1
X_16496_ _08968_ _09104_ vssd1 vssd1 vccd1 vccd1 _09106_ sky130_fd_sc_hd__nand2_1
XFILLER_206_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18235_ _02009_ _02010_ _02008_ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15447_ _07542_ _07592_ vssd1 vssd1 vccd1 vccd1 _08061_ sky130_fd_sc_hd__or2_1
X_12659_ _05310_ _05322_ _05329_ _05347_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__and4_1
XFILLER_54_1281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18166_ _01863_ _01864_ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__and2b_1
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15378_ _07509_ _07633_ _07991_ vssd1 vssd1 vccd1 vccd1 _07992_ sky130_fd_sc_hd__or3_1
XFILLER_157_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17117_ _09653_ _09655_ vssd1 vssd1 vccd1 vccd1 _09657_ sky130_fd_sc_hd__or2_1
X_14329_ _05431_ _07017_ vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__and2_1
XFILLER_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18097_ _01876_ _01877_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17048_ _09568_ _09588_ vssd1 vssd1 vccd1 vccd1 _09589_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18999_ rbzero.pov.spi_buffer\[47\] rbzero.pov.ready_buffer\[47\] _02651_ vssd1 vssd1
+ vccd1 vccd1 _02660_ sky130_fd_sc_hd__mux2_1
XFILLER_135_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20961_ net91 _00977_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20892_ net62 _00908_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_226_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21375_ _00398_ _01391_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20326_ _09247_ _03261_ _03262_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__and3_1
XFILLER_162_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20257_ _03254_ vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__clkinv_2
XFILLER_235_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20188_ rbzero.traced_texa\[3\] rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1 _03211_
+ sky130_fd_sc_hd__or2_1
XFILLER_114_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ net20 net19 _04670_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__and3_1
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13700_ _06388_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__clkbuf_4
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10912_ rbzero.tex_b0\[42\] rbzero.tex_b0\[41\] _03682_ vssd1 vssd1 vccd1 vccd1 _03683_
+ sky130_fd_sc_hd__mux2_1
XFILLER_245_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14680_ rbzero.wall_tracer.stepDistX\[-5\] _07185_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _07314_ sky130_fd_sc_hd__mux2_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11892_ rbzero.row_render.texu\[1\] _03289_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__or2_1
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13631_ _06260_ _06289_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__xor2_4
X_10843_ _03646_ vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13562_ _05866_ _06207_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__nor2_1
X_16350_ _08960_ _07537_ _07343_ vssd1 vssd1 vccd1 vccd1 _08961_ sky130_fd_sc_hd__mux2_1
XFILLER_125_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10774_ _03610_ vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15301_ _04937_ _07914_ vssd1 vssd1 vccd1 vccd1 _07915_ sky130_fd_sc_hd__or2_1
XFILLER_160_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12513_ _05146_ _05177_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__nor2_2
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16281_ _08889_ _08891_ vssd1 vssd1 vccd1 vccd1 _08892_ sky130_fd_sc_hd__and2_1
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13493_ _05401_ _05738_ _05854_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__and3_1
XFILLER_199_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18020_ _01682_ _01651_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__or2b_1
XFILLER_200_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15232_ _07836_ _07839_ _07844_ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__a21o_1
XFILLER_139_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12444_ _05133_ _05134_ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15163_ _07776_ _07745_ vssd1 vssd1 vccd1 vccd1 _07777_ sky130_fd_sc_hd__xnor2_1
XFILLER_166_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12375_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[11\] vssd1
+ vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__or2_1
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14114_ _06266_ _06634_ _06745_ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__o21bai_1
X_11326_ rbzero.row_render.size\[5\] rbzero.row_render.size\[4\] _04044_ vssd1 vssd1
+ vccd1 vccd1 _04045_ sky130_fd_sc_hd__or3_1
X_15094_ _07408_ _07702_ _07704_ _07707_ _04935_ vssd1 vssd1 vccd1 vccd1 _07708_ sky130_fd_sc_hd__a221o_1
XFILLER_141_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19971_ _03120_ vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__clkinv_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14045_ _06028_ _06305_ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__and2_1
XFILLER_119_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18922_ rbzero.pov.spi_buffer\[10\] rbzero.pov.ready_buffer\[10\] _02618_ vssd1 vssd1
+ vccd1 vccd1 _02620_ sky130_fd_sc_hd__mux2_1
X_11257_ rbzero.tex_r0\[37\] rbzero.tex_r0\[36\] _03974_ vssd1 vssd1 vccd1 vccd1 _03976_
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10208_ _03299_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__clkbuf_4
X_18853_ _02287_ _02565_ _02566_ _02569_ vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__a31o_1
XTAP_6460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11188_ _03853_ _03859_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__nand2_1
XTAP_6471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17804_ _10111_ _01587_ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__xor2_4
XTAP_6482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18784_ _02472_ rbzero.wall_tracer.rayAddendY\[5\] vssd1 vssd1 vccd1 vccd1 _02506_
+ sky130_fd_sc_hd__or2_1
XFILLER_209_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15996_ _08607_ _08608_ vssd1 vssd1 vccd1 vccd1 _08609_ sky130_fd_sc_hd__nor2_1
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17735_ _01424_ _01427_ _01517_ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__nand3_1
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14947_ rbzero.wall_tracer.visualWallDist\[-1\] _03795_ _07466_ vssd1 vssd1 vccd1
+ vccd1 _07561_ sky130_fd_sc_hd__a21oi_1
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17666_ _10116_ _10118_ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__nand2_1
XFILLER_165_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14878_ rbzero.debug_overlay.playerX\[-3\] _07411_ vssd1 vssd1 vccd1 vccd1 _07492_
+ sky130_fd_sc_hd__or2_1
XFILLER_90_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19405_ _02868_ vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__clkbuf_1
X_16617_ _09120_ _09225_ vssd1 vssd1 vccd1 vccd1 _09226_ sky130_fd_sc_hd__xnor2_1
XFILLER_211_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13829_ _06516_ _06517_ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__nand2_1
XFILLER_91_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17597_ _10001_ _10003_ vssd1 vssd1 vccd1 vccd1 _10134_ sky130_fd_sc_hd__nor2_1
XFILLER_23_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19336_ _02856_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__clkinv_2
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16548_ _09122_ _09123_ _09155_ vssd1 vssd1 vccd1 vccd1 _09157_ sky130_fd_sc_hd__nand3_1
XFILLER_143_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19267_ rbzero.spi_registers.new_other\[4\] rbzero.spi_registers.spi_buffer\[4\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__mux2_1
XFILLER_108_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16479_ _08974_ _09087_ _09088_ vssd1 vssd1 vccd1 vccd1 _09089_ sky130_fd_sc_hd__and3_1
XFILLER_223_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18218_ _05121_ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__clkbuf_4
XFILLER_178_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19198_ rbzero.spi_registers.vshift\[2\] _02774_ _02778_ _02738_ vssd1 vssd1 vccd1
+ vccd1 _00763_ sky130_fd_sc_hd__o211a_1
XFILLER_102_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18149_ _01857_ _01860_ _01858_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__o21a_1
XFILLER_129_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21160_ _00209_ _01176_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20111_ _03143_ _03146_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21091_ _00140_ _01107_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20042_ _03127_ vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__clkinv_2
XFILLER_59_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20944_ net76 _00960_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-9\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20875_ net58 _00891_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10490_ _03461_ vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12160_ _04853_ _04866_ _04860_ _04830_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__o211a_1
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21358_ _00381_ _01374_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ rbzero.traced_texVinit\[7\] rbzero.spi_registers.vshift\[4\] vssd1 vssd1
+ vccd1 vccd1 _03830_ sky130_fd_sc_hd__and2_1
X_20309_ rbzero.traced_texVinit\[0\] _09255_ _08573_ _09269_ vssd1 vssd1 vccd1 vccd1
+ _01394_ sky130_fd_sc_hd__o2bb2ai_1
X_12091_ _04789_ _04768_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__nor2_1
X_21289_ net114 _01305_ vssd1 vssd1 vccd1 vccd1 gpout5.clk_div\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ rbzero.otherx\[2\] _03736_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__xor2_1
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15850_ _07672_ _07673_ _07711_ _07400_ _07379_ vssd1 vssd1 vccd1 vccd1 _08464_ sky130_fd_sc_hd__a2111o_1
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _04936_ _07414_ vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__nand2_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15781_ _07645_ _08059_ _08393_ vssd1 vssd1 vccd1 vccd1 _08395_ sky130_fd_sc_hd__or3b_1
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12993_ _05678_ _05680_ _05681_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__nand3_1
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ _10056_ _08717_ _09920_ vssd1 vssd1 vccd1 vccd1 _10057_ sky130_fd_sc_hd__o21ba_1
XFILLER_206_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14732_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__buf_2
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11944_ net9 _04618_ net52 vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__and3_1
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _09733_ _09735_ _09988_ vssd1 vssd1 vccd1 vccd1 _09989_ sky130_fd_sc_hd__a21o_1
XFILLER_205_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14663_ _03800_ _07304_ _07305_ _07257_ vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__o211a_1
X_11875_ _04587_ _04588_ _04099_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__mux2_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16402_ _09010_ _09011_ vssd1 vssd1 vccd1 vccd1 _09012_ sky130_fd_sc_hd__nand2_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13614_ _06290_ _06288_ _06300_ _06302_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__a211oi_2
X_10826_ _03637_ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17382_ rbzero.wall_tracer.visualWallDist\[7\] _03796_ _08123_ vssd1 vssd1 vccd1
+ vccd1 _09920_ sky130_fd_sc_hd__and3_1
XFILLER_232_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14594_ rbzero.wall_tracer.visualWallDist\[-11\] _07253_ _07255_ _07256_ _07257_
+ vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__o221a_1
XFILLER_186_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19121_ rbzero.otherx\[2\] _02723_ _02730_ _02728_ vssd1 vssd1 vccd1 vccd1 _00734_
+ sky130_fd_sc_hd__o211a_1
X_16333_ _08941_ _08943_ vssd1 vssd1 vccd1 vccd1 _08944_ sky130_fd_sc_hd__xor2_1
XFILLER_186_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13545_ _06186_ _06187_ _06233_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__o21a_1
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10757_ rbzero.tex_g0\[51\] rbzero.tex_g0\[50\] _03593_ vssd1 vssd1 vccd1 vccd1 _03601_
+ sky130_fd_sc_hd__mux2_1
XFILLER_199_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19052_ _02687_ vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16264_ _08871_ _08873_ vssd1 vssd1 vccd1 vccd1 _08875_ sky130_fd_sc_hd__and2_1
X_13476_ _05936_ _06164_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__xor2_1
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10688_ _03565_ vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18003_ _10095_ _08735_ _01784_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__or3_1
XFILLER_200_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15215_ _07825_ _07828_ vssd1 vssd1 vccd1 vccd1 _07829_ sky130_fd_sc_hd__nand2_1
X_12427_ _05119_ rbzero.map_rom.c6 _05028_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__mux2_1
X_16195_ _08650_ _08651_ vssd1 vssd1 vccd1 vccd1 _08807_ sky130_fd_sc_hd__nor2_1
XFILLER_127_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15146_ _03795_ _07670_ _07466_ vssd1 vssd1 vccd1 vccd1 _07760_ sky130_fd_sc_hd__a21o_2
X_12358_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] rbzero.wall_tracer.rayAddendY\[5\]
+ rbzero.debug_overlay.facingY\[-3\] vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__o211a_1
XFILLER_181_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11309_ _03896_ _03955_ _03986_ _04006_ _04027_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__o32a_1
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15077_ _07689_ _07690_ vssd1 vssd1 vccd1 vccd1 _07691_ sky130_fd_sc_hd__nor2_1
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19954_ _03118_ vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__clkinv_2
X_12289_ _04951_ _04955_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__nand2_1
XFILLER_84_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14028_ _06516_ _06670_ _06668_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__nand3_1
X_18905_ rbzero.pov.spi_buffer\[2\] rbzero.pov.ready_buffer\[2\] _02608_ vssd1 vssd1
+ vccd1 vccd1 _02611_ sky130_fd_sc_hd__mux2_1
XFILLER_218_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19885_ _03111_ vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__clkinv_2
XFILLER_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18836_ rbzero.wall_tracer.rayAddendY\[8\] _00013_ _02554_ vssd1 vssd1 vccd1 vccd1
+ _00625_ sky130_fd_sc_hd__o21ba_1
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18767_ _02488_ _02489_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__nor2_1
XFILLER_209_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15979_ _08256_ vssd1 vssd1 vccd1 vccd1 _08592_ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17718_ _10023_ _10024_ _01501_ _01502_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__a31oi_1
XFILLER_209_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18698_ rbzero.wall_tracer.rayAddendY\[-1\] _02197_ _02425_ _02157_ vssd1 vssd1 vccd1
+ vccd1 _02426_ sky130_fd_sc_hd__a22o_1
XFILLER_236_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17649_ _01432_ _01433_ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__nand2_1
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20660_ net67 _00676_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_189_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19319_ _02849_ _02838_ _02850_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__and3b_1
XFILLER_52_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20591_ net96 _00607_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f4 sky130_fd_sc_hd__dfxtp_2
XFILLER_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21212_ _00261_ _01228_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21143_ _00192_ _01159_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21074_ _00123_ _01090_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20025_ _04702_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__buf_4
XFILLER_115_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20927_ net75 _00943_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[64\] sky130_fd_sc_hd__dfxtp_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11660_ rbzero.tex_g1\[25\] rbzero.tex_g1\[24\] _04374_ vssd1 vssd1 vccd1 vccd1 _04376_
+ sky130_fd_sc_hd__mux2_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20858_ _00076_ _00874_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[59\] sky130_fd_sc_hd__dfxtp_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10611_ rbzero.tex_g1\[56\] rbzero.tex_g1\[57\] _03519_ vssd1 vssd1 vccd1 vccd1 _03525_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11591_ _04306_ _04307_ _03909_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__mux2_1
XFILLER_168_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20789_ net101 _00805_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13330_ _05995_ _06017_ _06018_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__a21boi_1
XFILLER_126_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10542_ _03488_ vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13261_ _05949_ _05927_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ _03452_ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15000_ _07604_ _07612_ _07613_ vssd1 vssd1 vccd1 vccd1 _07614_ sky130_fd_sc_hd__a21o_1
XFILLER_170_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12212_ _04873_ _04883_ net38 net37 vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__or4_1
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13192_ _05839_ _05880_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__nor2_1
XFILLER_159_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12143_ net48 _04825_ _04820_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__and3_1
XFILLER_159_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16951_ _09423_ _09492_ vssd1 vssd1 vccd1 vccd1 _09493_ sky130_fd_sc_hd__xnor2_1
X_12074_ _04078_ _03781_ _03784_ _03291_ net21 _04773_ vssd1 vssd1 vccd1 vccd1 _04782_
+ sky130_fd_sc_hd__mux4_1
XFILLER_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15902_ _07388_ _07567_ vssd1 vssd1 vccd1 vccd1 _08516_ sky130_fd_sc_hd__or2_1
X_11025_ _03736_ rbzero.map_rom.f1 _03752_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__or3_1
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19670_ _02727_ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__buf_4
XFILLER_46_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16882_ _09174_ _09175_ vssd1 vssd1 vccd1 vccd1 _09424_ sky130_fd_sc_hd__nor2_1
XFILLER_77_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18621_ _02353_ _02354_ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__nand2_1
XFILLER_77_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15833_ _08353_ _08354_ _08446_ vssd1 vssd1 vccd1 vccd1 _08447_ sky130_fd_sc_hd__a21o_1
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18552_ _02293_ _02294_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__nand2_1
X_15764_ _08288_ _08376_ vssd1 vssd1 vccd1 vccd1 _08378_ sky130_fd_sc_hd__and2b_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _05656_ _05664_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__xnor2_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17503_ _08507_ _09115_ _09915_ _09916_ vssd1 vssd1 vccd1 vccd1 _10040_ sky130_fd_sc_hd__o31a_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _04940_ vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__buf_4
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _04623_ _04627_ _04637_ net11 vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__a22o_1
X_18483_ _09261_ _02221_ _02222_ _02230_ vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__a31o_1
X_15695_ _08287_ _08308_ vssd1 vssd1 vccd1 vccd1 _08309_ sky130_fd_sc_hd__xor2_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _09954_ _09971_ vssd1 vssd1 vccd1 vccd1 _09972_ sky130_fd_sc_hd__xor2_1
XFILLER_221_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14646_ rbzero.wall_tracer.trackDistX\[5\] vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__inv_2
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ _04570_ _04571_ _03915_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__mux2_1
XFILLER_53_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17365_ _09796_ _09806_ _09804_ vssd1 vssd1 vccd1 vccd1 _09903_ sky130_fd_sc_hd__a21o_1
XFILLER_202_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10809_ rbzero.tex_g0\[27\] rbzero.tex_g0\[26\] _03627_ vssd1 vssd1 vccd1 vccd1 _03629_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_19 rbzero.pov.mosi vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14577_ _05440_ _07007_ _07038_ _07101_ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__and4_1
XFILLER_14_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11789_ rbzero.tex_b0\[7\] _04143_ _04145_ _03930_ vssd1 vssd1 vccd1 vccd1 _04504_
+ sky130_fd_sc_hd__a31o_1
XFILLER_159_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19104_ gpout0.vpos\[2\] gpout0.vpos\[1\] gpout0.vpos\[0\] vssd1 vssd1 vccd1 vccd1
+ _02716_ sky130_fd_sc_hd__and3_1
X_16316_ _08915_ _08926_ vssd1 vssd1 vccd1 vccd1 _08927_ sky130_fd_sc_hd__xnor2_1
XFILLER_192_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13528_ _06178_ _06216_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__xor2_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17296_ _09832_ _09834_ vssd1 vssd1 vccd1 vccd1 _09835_ sky130_fd_sc_hd__xnor2_1
XFILLER_185_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19035_ rbzero.pov.spi_buffer\[64\] rbzero.pov.ready_buffer\[64\] _02673_ vssd1 vssd1
+ vccd1 vccd1 _02679_ sky130_fd_sc_hd__mux2_1
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16247_ _08429_ _08724_ vssd1 vssd1 vccd1 vccd1 _08858_ sky130_fd_sc_hd__or2_1
XFILLER_173_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13459_ _06066_ _06067_ _06147_ _06095_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__and4bb_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16178_ _08779_ _08636_ _08786_ _08789_ vssd1 vssd1 vccd1 vccd1 _08790_ sky130_fd_sc_hd__nand4_1
XFILLER_115_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15129_ _07742_ _07400_ vssd1 vssd1 vccd1 vccd1 _07743_ sky130_fd_sc_hd__nor2_1
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19937_ _03114_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__buf_4
XFILLER_190_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19868_ _03109_ vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__clkinv_2
XFILLER_233_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18819_ _02537_ _02538_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__nand2_1
XFILLER_56_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19799_ gpout0.vpos\[7\] gpout0.vpos\[6\] _03096_ vssd1 vssd1 vccd1 vccd1 _03099_
+ sky130_fd_sc_hd__and3_1
XFILLER_243_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20712_ net99 _00728_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.ss_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20643_ net66 _00659_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20574_ net89 _00590_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21126_ _00175_ _01142_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21057_ _00106_ _01073_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20008_ _03123_ vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__clkinv_2
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12830_ _05517_ _05451_ _05518_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__a21boi_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _05333_ _05334_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__or2_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _05527_ _07151_ _07177_ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__a21o_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ rbzero.tex_g1\[47\] _03964_ _03965_ _03997_ vssd1 vssd1 vccd1 vccd1 _04428_
+ sky130_fd_sc_hd__a31o_1
XFILLER_230_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15480_ _08050_ _08051_ vssd1 vssd1 vccd1 vccd1 _08094_ sky130_fd_sc_hd__xnor2_1
X_12692_ _05260_ _05380_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__xnor2_4
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _07119_ vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__clkbuf_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _03972_ _04355_ _04359_ _03950_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__a211o_1
XFILLER_74_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17150_ _09678_ _09689_ vssd1 vssd1 vccd1 vccd1 _09690_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14362_ _05408_ _07050_ vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__or2_1
XFILLER_168_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11574_ rbzero.debug_overlay.playerX\[3\] _04231_ _04209_ rbzero.debug_overlay.playerX\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__a22o_1
XFILLER_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput17 i_gpout2_sel[2] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_6
X_16101_ _08680_ _08681_ _08712_ vssd1 vssd1 vccd1 vccd1 _08713_ sky130_fd_sc_hd__o21ai_1
XFILLER_183_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput28 i_gpout4_sel[1] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_6
XFILLER_156_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13313_ _05627_ _05616_ _05657_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__or3_2
X_10525_ rbzero.tex_r0\[34\] rbzero.tex_r0\[33\] _03479_ vssd1 vssd1 vccd1 vccd1 _03480_
+ sky130_fd_sc_hd__mux2_1
Xinput39 i_mode[0] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_6
X_17081_ _09619_ _09621_ vssd1 vssd1 vccd1 vccd1 _09622_ sky130_fd_sc_hd__xnor2_1
X_14293_ _06455_ _06974_ _06453_ vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__a21boi_1
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16032_ _08644_ vssd1 vssd1 vccd1 vccd1 _08645_ sky130_fd_sc_hd__buf_4
X_13244_ _05834_ _05836_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__xor2_1
XFILLER_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10456_ _03441_ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13175_ _05692_ _05710_ _05772_ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__a31oi_1
XFILLER_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10387_ _03405_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12126_ _04078_ _03781_ _03784_ _03291_ net27 _04825_ vssd1 vssd1 vccd1 vccd1 _04833_
+ sky130_fd_sc_hd__mux4_1
XFILLER_170_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17983_ _08123_ _09115_ vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__nor2_1
XFILLER_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19722_ rbzero.pov.ready_buffer\[42\] _03056_ _03059_ rbzero.debug_overlay.facingX\[0\]
+ _03065_ vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__o221a_1
X_16934_ _09201_ _09474_ _09475_ vssd1 vssd1 vccd1 vccd1 _09476_ sky130_fd_sc_hd__and3_1
X_12057_ net5 _04735_ _04758_ _04765_ _04753_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__a32o_1
XFILLER_81_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11008_ rbzero.map_rom.f2 vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__clkbuf_4
XFILLER_77_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19653_ _07360_ _02958_ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__nor2_1
XFILLER_77_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16865_ _08086_ _08223_ _07620_ _08671_ vssd1 vssd1 vccd1 vccd1 _09407_ sky130_fd_sc_hd__or4_1
XFILLER_133_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18604_ _02337_ _02325_ _02329_ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__and3b_1
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15816_ _07625_ _07680_ _07847_ _08429_ vssd1 vssd1 vccd1 vccd1 _08430_ sky130_fd_sc_hd__o22a_1
X_19584_ rbzero.pov.ready_buffer\[61\] _07464_ _02963_ vssd1 vssd1 vccd1 vccd1 _02966_
+ sky130_fd_sc_hd__mux2_1
X_16796_ _09332_ _09334_ _09333_ vssd1 vssd1 vccd1 vccd1 _09342_ sky130_fd_sc_hd__a21boi_1
XFILLER_203_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18535_ _02277_ _02278_ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__nand2_1
XFILLER_234_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15747_ _07435_ _08296_ _07971_ _07986_ vssd1 vssd1 vccd1 vccd1 _08361_ sky130_fd_sc_hd__or4_1
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _05645_ _05634_ _05646_ _05647_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__a31o_1
XFILLER_46_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18466_ _02208_ _02213_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__nand2_1
XFILLER_233_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15678_ _08255_ _08257_ vssd1 vssd1 vccd1 vccd1 _08292_ sky130_fd_sc_hd__xnor2_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17417_ _07663_ vssd1 vssd1 vccd1 vccd1 _09955_ sky130_fd_sc_hd__clkbuf_4
X_14629_ rbzero.wall_tracer.trackDistX\[0\] rbzero.wall_tracer.trackDistY\[0\] _07258_
+ vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__mux2_1
XFILLER_18_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18397_ _02147_ _02150_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__and2_1
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17348_ _09885_ _09886_ vssd1 vssd1 vccd1 vccd1 _09887_ sky130_fd_sc_hd__xnor2_4
XFILLER_202_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17279_ _09808_ _09817_ vssd1 vssd1 vccd1 vccd1 _09818_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19018_ rbzero.pov.spi_buffer\[56\] rbzero.pov.ready_buffer\[56\] _02662_ vssd1 vssd1
+ vccd1 vccd1 _02670_ sky130_fd_sc_hd__mux2_1
XFILLER_106_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20290_ _03257_ vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__clkinv_2
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20626_ net54 _00642_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20557_ net123 _00573_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10310_ _03364_ vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11290_ rbzero.tex_r0\[13\] rbzero.tex_r0\[12\] _03961_ vssd1 vssd1 vccd1 vccd1 _04009_
+ sky130_fd_sc_hd__mux2_1
X_20488_ net112 _00504_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10241_ _03328_ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21109_ _00158_ _01125_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_6867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14980_ _07591_ _07593_ vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__nor2_1
XTAP_6889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13931_ _06604_ _06619_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16650_ _09250_ vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__clkbuf_1
X_13862_ _05434_ _06550_ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__nor2_1
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15601_ _08189_ _08214_ vssd1 vssd1 vccd1 vccd1 _08215_ sky130_fd_sc_hd__xor2_2
XFILLER_170_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12813_ _05395_ _05378_ _05429_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__mux2_1
X_16581_ _07824_ _08793_ _08272_ vssd1 vssd1 vccd1 vccd1 _09190_ sky130_fd_sc_hd__a21oi_1
XFILLER_216_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13793_ _06174_ _06481_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__nor2_1
XFILLER_215_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18320_ _02082_ _02083_ _02084_ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__and3_1
XFILLER_43_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15532_ _08131_ _08144_ vssd1 vssd1 vccd1 vccd1 _08146_ sky130_fd_sc_hd__and2b_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12744_ _05336_ _05416_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__nor2_2
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18251_ _01997_ _02024_ _02025_ _02013_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__a31o_1
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _08021_ _08019_ _08020_ vssd1 vssd1 vccd1 vccd1 _08077_ sky130_fd_sc_hd__a21oi_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _05237_ _05239_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__and2_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17202_ _09601_ _09618_ _09741_ vssd1 vssd1 vccd1 vccd1 _09742_ sky130_fd_sc_hd__a21bo_1
X_14414_ _06997_ _06994_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__or2_1
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18182_ _01945_ _01961_ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__xnor2_1
XFILLER_198_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11626_ _04339_ _04342_ _03923_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__mux2_1
X_15394_ _07350_ _07353_ _07354_ _07644_ vssd1 vssd1 vccd1 vccd1 _08008_ sky130_fd_sc_hd__a211o_1
XFILLER_54_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17133_ _08599_ _08725_ _09538_ _09537_ vssd1 vssd1 vccd1 vccd1 _09673_ sky130_fd_sc_hd__o31a_1
XFILLER_15_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14345_ _06981_ _06996_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__and2_1
XFILLER_128_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11557_ gpout0.vpos\[3\] _04252_ _04259_ _04267_ _04274_ vssd1 vssd1 vccd1 vccd1
+ _04275_ sky130_fd_sc_hd__a221o_1
XFILLER_7_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17064_ _07814_ _09463_ _09467_ _09603_ vssd1 vssd1 vccd1 vccd1 _09605_ sky130_fd_sc_hd__o22ai_1
X_10508_ rbzero.tex_r0\[42\] rbzero.tex_r0\[41\] _03468_ vssd1 vssd1 vccd1 vccd1 _03471_
+ sky130_fd_sc_hd__mux2_1
X_14276_ _06790_ _06782_ _06788_ vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__and3_1
X_11488_ _03293_ _04205_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__nand2_2
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16015_ _07663_ _08484_ vssd1 vssd1 vccd1 vccd1 _08628_ sky130_fd_sc_hd__and2_2
X_13227_ _05796_ _05911_ _05912_ _05915_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__a2bb2o_1
X_10439_ _03432_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13158_ _05645_ _05567_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__and2_1
XFILLER_112_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12109_ _04785_ net23 _04813_ _04816_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__a31o_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17966_ _01746_ _01747_ vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__xor2_1
X_13089_ _05765_ _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16917_ _09457_ _09458_ vssd1 vssd1 vccd1 vccd1 _09459_ sky130_fd_sc_hd__and2_1
X_19705_ _03058_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__buf_2
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17897_ _01548_ _01555_ _01679_ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__a21oi_1
XFILLER_211_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16848_ _08429_ _09389_ vssd1 vssd1 vccd1 vccd1 _09390_ sky130_fd_sc_hd__nand2_1
X_19636_ rbzero.pov.ready_buffer\[73\] _02836_ _02955_ _03005_ vssd1 vssd1 vccd1 vccd1
+ _03006_ sky130_fd_sc_hd__a211o_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19567_ _02952_ vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__clkbuf_1
XFILLER_241_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16779_ _09318_ _09320_ _09319_ vssd1 vssd1 vccd1 vccd1 _09327_ sky130_fd_sc_hd__a21boi_1
XFILLER_111_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18518_ _02191_ rbzero.debug_overlay.vplaneX\[-5\] _02261_ _02262_ vssd1 vssd1 vccd1
+ vccd1 _02263_ sky130_fd_sc_hd__o22ai_1
XFILLER_55_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19498_ rbzero.pov.spi_buffer\[45\] rbzero.pov.spi_buffer\[46\] _02910_ vssd1 vssd1
+ vccd1 vccd1 _02917_ sky130_fd_sc_hd__mux2_1
XFILLER_185_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18449_ rbzero.debug_overlay.vplaneX\[-5\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__nand2_1
XFILLER_178_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20411_ net130 _00442_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_21391_ net110 _01407_ vssd1 vssd1 vccd1 vccd1 gpout0.clk_div\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20342_ rbzero.wall_tracer.rayAddendX\[-6\] _03260_ _09267_ _03272_ vssd1 vssd1 vccd1
+ vccd1 _01413_ sky130_fd_sc_hd__a22o_1
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20273_ _03256_ vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__clkinv_2
XFILLER_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10790_ rbzero.tex_g0\[36\] rbzero.tex_g0\[35\] _03616_ vssd1 vssd1 vccd1 vccd1 _03619_
+ sky130_fd_sc_hd__mux2_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12460_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__nand2_2
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11411_ _04127_ _04128_ _03942_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__mux2_1
XFILLER_197_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12391_ _05075_ _05083_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__and2_1
X_20609_ net90 _00625_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14130_ _06764_ _06818_ vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__xor2_1
XFILLER_181_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11342_ _04055_ gpout0.hpos\[3\] gpout0.hpos\[4\] _04054_ _04060_ vssd1 vssd1 vccd1
+ vccd1 _04061_ sky130_fd_sc_hd__a221o_1
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14061_ _06636_ _06749_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__or2_1
X_11273_ _03990_ _03991_ _03957_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__mux2_1
XFILLER_153_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13012_ _05700_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__buf_2
X_10224_ _03319_ vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17820_ _10161_ _01493_ _01491_ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__a21oi_1
XTAP_6642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17751_ _07472_ _08663_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__or2_1
XFILLER_121_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14963_ _07556_ _07576_ vssd1 vssd1 vccd1 vccd1 _07577_ sky130_fd_sc_hd__xnor2_1
XTAP_5974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16702_ rbzero.traced_texa\[4\] _09264_ _09265_ rbzero.wall_tracer.visualWallDist\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__a22o_1
XFILLER_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13914_ _06532_ _06533_ _06534_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__o21ai_1
X_17682_ _01464_ _01466_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__xor2_1
XFILLER_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14894_ _07507_ vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__buf_2
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19421_ _02876_ vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__clkbuf_1
X_16633_ rbzero.wall_tracer.texu\[5\] _07338_ vssd1 vssd1 vccd1 vccd1 _09242_ sky130_fd_sc_hd__or2_1
XFILLER_223_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13845_ _06520_ _06519_ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__xor2_1
XFILLER_235_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19352_ _02858_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__clkinv_2
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16564_ _07751_ _07834_ _09170_ _09171_ _09172_ vssd1 vssd1 vccd1 vccd1 _09173_ sky130_fd_sc_hd__o32a_1
XFILLER_188_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13776_ _06462_ _06463_ _06464_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__nand3_1
XFILLER_203_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10988_ _03722_ vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__clkbuf_1
XFILLER_206_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18303_ rbzero.wall_tracer.trackDistY\[0\] rbzero.wall_tracer.stepDistY\[0\] vssd1
+ vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__or2_1
X_15515_ _08126_ _08128_ vssd1 vssd1 vccd1 vccd1 _08129_ sky130_fd_sc_hd__xor2_1
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12727_ _05361_ _05363_ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__or2_2
X_19283_ _02826_ vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16495_ _08968_ _09104_ vssd1 vssd1 vccd1 vccd1 _09105_ sky130_fd_sc_hd__or2_1
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18234_ _02008_ _02009_ _02010_ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__or3_1
X_15446_ _08059_ vssd1 vssd1 vccd1 vccd1 _08060_ sky130_fd_sc_hd__buf_2
XFILLER_129_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12658_ _05335_ _05344_ _05346_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__and3b_1
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18165_ _01941_ _01944_ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__xnor2_1
X_11609_ rbzero.tex_g0\[7\] _03939_ _03941_ _04014_ vssd1 vssd1 vccd1 vccd1 _04326_
+ sky130_fd_sc_hd__a31o_1
XFILLER_102_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15377_ _07501_ _07986_ vssd1 vssd1 vccd1 vccd1 _07991_ sky130_fd_sc_hd__or2_1
X_12589_ rbzero.wall_tracer.visualWallDist\[7\] _05190_ vssd1 vssd1 vccd1 vccd1 _05278_
+ sky130_fd_sc_hd__and2_1
XFILLER_128_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17116_ _09653_ _09655_ vssd1 vssd1 vccd1 vccd1 _09656_ sky130_fd_sc_hd__nand2_1
XFILLER_184_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14328_ _06690_ _06970_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__xor2_1
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18096_ _07827_ _07914_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__nor2_1
XFILLER_209_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17047_ _09586_ _09587_ vssd1 vssd1 vccd1 vccd1 _09588_ sky130_fd_sc_hd__or2b_1
XFILLER_132_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14259_ _06844_ _06914_ _06920_ _06947_ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__o211a_1
XFILLER_217_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18998_ _02659_ vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__clkbuf_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17949_ _01591_ _01621_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__and2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20960_ net91 _00976_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_226_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19619_ _02990_ _02835_ _02991_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__or3b_1
XFILLER_226_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20891_ net64 _00907_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_246_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21374_ _00397_ _01390_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20325_ gpout0.clk_div\[0\] gpout0.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__or2_1
XFILLER_235_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20256_ _03254_ vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__clkinv_2
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20187_ _09245_ _03208_ _03210_ _03064_ rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1
+ _01320_ sky130_fd_sc_hd__a32o_1
XTAP_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ net16 net17 net18 vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__a21o_1
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ _03604_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__clkbuf_4
XFILLER_232_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ _04591_ _04592_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__nor2_1
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13630_ _06317_ _06318_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__or2_1
XFILLER_232_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10842_ rbzero.tex_g0\[11\] rbzero.tex_g0\[10\] _03638_ vssd1 vssd1 vccd1 vccd1 _03646_
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13561_ _06229_ _06249_ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10773_ rbzero.tex_g0\[44\] rbzero.tex_g0\[43\] _03605_ vssd1 vssd1 vccd1 vccd1 _03610_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15300_ rbzero.wall_tracer.visualWallDist\[5\] _03795_ vssd1 vssd1 vccd1 vccd1 _07914_
+ sky130_fd_sc_hd__nand2_4
XFILLER_164_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12512_ rbzero.wall_tracer.visualWallDist\[1\] _05190_ _03789_ vssd1 vssd1 vccd1
+ vccd1 _05201_ sky130_fd_sc_hd__a21oi_2
X_16280_ _08890_ _07886_ _08888_ vssd1 vssd1 vccd1 vccd1 _08891_ sky130_fd_sc_hd__o21ai_1
XFILLER_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13492_ _05756_ _05855_ _06180_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__a21o_1
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15231_ _07836_ _07839_ _07844_ vssd1 vssd1 vccd1 vccd1 _07845_ sky130_fd_sc_hd__nand3_1
XFILLER_173_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12443_ _05122_ _05127_ vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__nand2_1
XFILLER_51_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15162_ _07380_ _07743_ _07744_ vssd1 vssd1 vccd1 vccd1 _07776_ sky130_fd_sc_hd__a21boi_1
XFILLER_154_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12374_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[11\] vssd1
+ vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__nand2_1
XFILLER_193_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14113_ _06798_ _06799_ _06800_ _06801_ vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__a22o_1
X_11325_ rbzero.row_render.size\[3\] _04043_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__or2_1
XFILLER_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15093_ _07351_ _07706_ vssd1 vssd1 vccd1 vccd1 _07707_ sky130_fd_sc_hd__nor2_1
XFILLER_153_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19970_ _03114_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__clkbuf_8
XFILLER_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14044_ _06706_ _06732_ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__xnor2_2
XFILLER_158_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11256_ rbzero.tex_r0\[39\] rbzero.tex_r0\[38\] _03974_ vssd1 vssd1 vccd1 vccd1 _03975_
+ sky130_fd_sc_hd__mux2_1
X_18921_ _02619_ vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__clkbuf_1
XTAP_7140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ _03310_ vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11187_ rbzero.tex_r0\[51\] rbzero.tex_r0\[50\] _03904_ vssd1 vssd1 vccd1 vccd1 _03906_
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18852_ rbzero.wall_tracer.rayAddendY\[10\] _02158_ _02568_ vssd1 vssd1 vccd1 vccd1
+ _02569_ sky130_fd_sc_hd__a21bo_1
XTAP_6450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17803_ _09182_ _01585_ _01586_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__mux2_2
XTAP_6483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18783_ _02472_ rbzero.wall_tracer.rayAddendY\[5\] vssd1 vssd1 vccd1 vccd1 _02505_
+ sky130_fd_sc_hd__nand2_1
X_15995_ _07388_ _07805_ _08515_ _08513_ vssd1 vssd1 vccd1 vccd1 _08608_ sky130_fd_sc_hd__o31a_1
XTAP_5760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17734_ _01424_ _01427_ _01517_ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__a21o_1
XTAP_5782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14946_ _07453_ _07559_ vssd1 vssd1 vccd1 vccd1 _07560_ sky130_fd_sc_hd__nand2_1
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17665_ _10099_ _10106_ _01449_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__a21o_1
XFILLER_208_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14877_ _07374_ vssd1 vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__buf_4
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16616_ _09223_ _09224_ vssd1 vssd1 vccd1 vccd1 _09225_ sky130_fd_sc_hd__xor2_1
X_19404_ rbzero.pov.spi_buffer\[0\] rbzero.pov.spi_buffer\[1\] _02866_ vssd1 vssd1
+ vccd1 vccd1 _02868_ sky130_fd_sc_hd__mux2_1
X_13828_ _06471_ _06472_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__xor2_1
X_17596_ _10090_ _10132_ vssd1 vssd1 vccd1 vccd1 _10133_ sky130_fd_sc_hd__xnor2_1
XFILLER_223_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16547_ _09122_ _09123_ _09155_ vssd1 vssd1 vccd1 vccd1 _09156_ sky130_fd_sc_hd__a21o_1
XFILLER_206_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19335_ _02856_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__clkinv_2
XFILLER_232_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13759_ _06446_ _06447_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__nor2_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19266_ _02817_ vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__clkbuf_1
X_16478_ _09083_ _09084_ _09086_ vssd1 vssd1 vccd1 vccd1 _09088_ sky130_fd_sc_hd__a21o_1
XFILLER_203_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18217_ _01995_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__clkbuf_4
X_15429_ _07967_ _07965_ vssd1 vssd1 vccd1 vccd1 _08043_ sky130_fd_sc_hd__and2b_1
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19197_ rbzero.spi_registers.new_vshift\[2\] _02775_ vssd1 vssd1 vccd1 vccd1 _02778_
+ sky130_fd_sc_hd__or2_1
XFILLER_223_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18148_ _08594_ _09976_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__nor2_1
XFILLER_8_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18079_ _09429_ _09389_ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__nand2_1
XFILLER_117_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20110_ _03144_ _03145_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__and2b_1
XFILLER_144_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21090_ _00139_ _01106_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20041_ _03127_ vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__clkinv_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20943_ net85 _00959_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20874_ net58 _00890_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21357_ _00380_ _01373_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11110_ rbzero.texV\[6\] _03827_ _03828_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__nand3_1
XFILLER_155_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20308_ _02855_ vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__clkinv_2
X_12090_ _04789_ net21 vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__and2_1
XFILLER_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21288_ net114 _01304_ vssd1 vssd1 vccd1 vccd1 gpout5.clk_div\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_235_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11041_ rbzero.othery\[1\] rbzero.map_rom.c6 vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__xor2_1
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20239_ _03125_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__buf_4
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ _07410_ _07413_ _07374_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__mux2_1
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15780_ _07646_ _08059_ _08393_ vssd1 vssd1 vccd1 vccd1 _08394_ sky130_fd_sc_hd__o21ba_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12992_ _05634_ _05636_ _05611_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__a21oi_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14731_ _07100_ _07187_ _07188_ _07336_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__a31o_1
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ _04115_ _04651_ _04653_ gpout1.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _04654_
+ sky130_fd_sc_hd__a22o_1
XFILLER_245_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _09987_ _07814_ _09857_ vssd1 vssd1 vccd1 vccd1 _09988_ sky130_fd_sc_hd__mux2_1
XFILLER_205_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14662_ _05301_ _03800_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__nand2_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11874_ rbzero.color_sky\[5\] rbzero.color_floor\[5\] _04030_ vssd1 vssd1 vccd1 vccd1
+ _04588_ sky130_fd_sc_hd__mux2_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _08976_ _08977_ _09009_ vssd1 vssd1 vccd1 vccd1 _09011_ sky130_fd_sc_hd__nand3_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13613_ _06287_ _06301_ _06285_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__a21o_1
XFILLER_72_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17381_ _09917_ _09918_ vssd1 vssd1 vccd1 vccd1 _09919_ sky130_fd_sc_hd__xnor2_1
X_10825_ rbzero.tex_g0\[19\] rbzero.tex_g0\[18\] _03627_ vssd1 vssd1 vccd1 vccd1 _03637_
+ sky130_fd_sc_hd__mux2_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14593_ _03819_ vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__clkbuf_4
XFILLER_60_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19120_ rbzero.spi_registers.new_other\[8\] _02725_ vssd1 vssd1 vccd1 vccd1 _02730_
+ sky130_fd_sc_hd__or2_1
X_16332_ _08778_ _08805_ _08942_ vssd1 vssd1 vccd1 vccd1 _08943_ sky130_fd_sc_hd__a21o_1
XFILLER_158_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13544_ _06231_ _06232_ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__and2_1
XFILLER_125_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10756_ _03600_ vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19051_ rbzero.pov.spi_buffer\[72\] rbzero.pov.ready_buffer\[72\] _02607_ vssd1 vssd1
+ vccd1 vccd1 _02687_ sky130_fd_sc_hd__mux2_1
X_16263_ _08871_ _08873_ vssd1 vssd1 vccd1 vccd1 _08874_ sky130_fd_sc_hd__nor2_1
XFILLER_125_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13475_ _05881_ _05980_ _06161_ _06163_ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__a22o_1
XFILLER_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10687_ rbzero.tex_g1\[20\] rbzero.tex_g1\[21\] _03563_ vssd1 vssd1 vccd1 vccd1 _03565_
+ sky130_fd_sc_hd__mux2_1
X_18002_ _01782_ _01783_ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__xnor2_1
X_15214_ _07826_ _07817_ _07827_ _07471_ vssd1 vssd1 vccd1 vccd1 _07828_ sky130_fd_sc_hd__o22ai_1
XFILLER_51_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12426_ rbzero.debug_overlay.playerY\[1\] _05118_ _03798_ vssd1 vssd1 vccd1 vccd1
+ _05119_ sky130_fd_sc_hd__mux2_1
XFILLER_127_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16194_ _08778_ _08805_ vssd1 vssd1 vccd1 vccd1 _08806_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15145_ _07645_ _07675_ _07708_ _07735_ vssd1 vssd1 vccd1 vccd1 _07759_ sky130_fd_sc_hd__or4_1
X_12357_ _05045_ _05049_ _05034_ _05033_ _05030_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__a2111oi_1
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11308_ _03985_ _04017_ _04025_ _04026_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__a31o_1
X_15076_ _07446_ _07448_ _07655_ _07656_ _07447_ vssd1 vssd1 vccd1 vccd1 _07690_ sky130_fd_sc_hd__o2111a_1
X_19953_ _03118_ vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__clkinv_2
X_12288_ _04975_ _04976_ _04978_ _04981_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__o31a_1
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14027_ _06715_ _06693_ vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__xnor2_1
X_18904_ _02610_ vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__clkbuf_1
XFILLER_214_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11239_ _03957_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__clkbuf_4
X_19884_ _03111_ vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__clkinv_2
XFILLER_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18835_ _03729_ _02546_ _02553_ _03812_ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__o211a_1
XTAP_6280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15978_ _08461_ _08470_ _08468_ vssd1 vssd1 vccd1 vccd1 _08591_ sky130_fd_sc_hd__a21o_1
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18766_ _02473_ _02478_ _02487_ _03729_ vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__a31o_1
XTAP_5590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17717_ _10018_ _10144_ _10143_ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__a21o_1
XFILLER_236_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14929_ rbzero.debug_overlay.playerY\[-2\] _07497_ vssd1 vssd1 vccd1 vccd1 _07543_
+ sky130_fd_sc_hd__xor2_1
XFILLER_247_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18697_ _02414_ _02424_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17648_ _07618_ _07663_ _10074_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__or3b_1
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17579_ _10111_ _10114_ _10115_ vssd1 vssd1 vccd1 vccd1 _10116_ sky130_fd_sc_hd__nand3_1
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19318_ rbzero.pov.spi_counter\[3\] rbzero.pov.spi_counter\[2\] _02840_ rbzero.pov.spi_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__a31o_1
XFILLER_143_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20590_ net95 _00606_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19249_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.new_leak\[3\] _02804_
+ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__mux2_1
XFILLER_108_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21211_ _00260_ _01227_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21142_ _00191_ _01158_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21073_ _00122_ _01089_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20024_ _03124_ vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__clkinv_2
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20926_ net75 _00942_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[63\] sky130_fd_sc_hd__dfxtp_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20857_ _00075_ _00873_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _03524_ vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_211_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11590_ rbzero.tex_g0\[23\] rbzero.tex_g0\[22\] _04119_ vssd1 vssd1 vccd1 vccd1 _04307_
+ sky130_fd_sc_hd__mux2_1
XFILLER_195_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20788_ net102 _00804_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10541_ rbzero.tex_r0\[26\] rbzero.tex_r0\[25\] _03479_ vssd1 vssd1 vccd1 vccd1 _03488_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13260_ _05906_ _05924_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__xnor2_1
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10472_ rbzero.tex_r0\[59\] rbzero.tex_r0\[58\] _03446_ vssd1 vssd1 vccd1 vccd1 _03452_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12211_ _04892_ _04894_ _04898_ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__a31o_1
X_13191_ _05838_ _05784_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__and2b_1
XFILLER_151_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12142_ _04840_ _04820_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__nor2_1
XFILLER_150_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16950_ _09489_ _09491_ vssd1 vssd1 vccd1 vccd1 _09492_ sky130_fd_sc_hd__xnor2_1
XFILLER_150_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12073_ net26 net25 _04780_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__and3_1
XFILLER_151_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15901_ _08513_ _08514_ vssd1 vssd1 vccd1 vccd1 _08515_ sky130_fd_sc_hd__nand2_1
XFILLER_172_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11024_ rbzero.map_rom.f4 rbzero.map_rom.f3 rbzero.map_rom.i_col\[4\] vssd1 vssd1
+ vccd1 vccd1 _03752_ sky130_fd_sc_hd__or3_1
XFILLER_81_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16881_ _09383_ _09422_ vssd1 vssd1 vccd1 vccd1 _09423_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15832_ _08271_ _08314_ vssd1 vssd1 vccd1 vccd1 _08446_ sky130_fd_sc_hd__nor2_1
X_18620_ _02353_ _02354_ vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__or2_1
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15763_ _08376_ _08288_ vssd1 vssd1 vccd1 vccd1 _08377_ sky130_fd_sc_hd__and2b_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ _02247_ rbzero.debug_overlay.vplaneX\[-3\] rbzero.debug_overlay.vplaneX\[-2\]
+ vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__or3b_1
X_12975_ _05658_ _05660_ _05661_ _05663_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__o22ai_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17502_ _09949_ _09913_ vssd1 vssd1 vccd1 vccd1 _10039_ sky130_fd_sc_hd__or2b_1
X_14714_ _07331_ vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__clkbuf_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ _04618_ net12 _04629_ _04634_ _04636_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__a32o_1
X_18482_ rbzero.wall_tracer.rayAddendX\[1\] _02197_ _02229_ _02157_ vssd1 vssd1 vccd1
+ vccd1 _02230_ sky130_fd_sc_hd__a22o_1
X_15694_ _08290_ _08306_ _08307_ vssd1 vssd1 vccd1 vccd1 _08308_ sky130_fd_sc_hd__a21boi_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _09960_ _09970_ vssd1 vssd1 vccd1 vccd1 _09971_ sky130_fd_sc_hd__xnor2_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _05002_ _07254_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__nor2_1
XFILLER_60_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ rbzero.tex_b1\[13\] rbzero.tex_b1\[12\] _04544_ vssd1 vssd1 vccd1 vccd1 _04571_
+ sky130_fd_sc_hd__mux2_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17364_ _09824_ _09789_ vssd1 vssd1 vccd1 vccd1 _09902_ sky130_fd_sc_hd__or2b_1
X_10808_ _03628_ vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14576_ _07242_ vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11788_ rbzero.tex_b0\[6\] _03959_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__and2_1
XFILLER_202_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16315_ _08924_ _08925_ vssd1 vssd1 vccd1 vccd1 _08926_ sky130_fd_sc_hd__nor2_1
XFILLER_14_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19103_ _02715_ vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__clkbuf_1
X_13527_ _06214_ _06215_ vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__nor2_1
XFILLER_140_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17295_ _09833_ _07631_ vssd1 vssd1 vccd1 vccd1 _09834_ sky130_fd_sc_hd__nor2_1
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10739_ _03591_ vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19034_ _02678_ vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__clkbuf_1
X_16246_ _08854_ _08856_ vssd1 vssd1 vccd1 vccd1 _08857_ sky130_fd_sc_hd__nand2_1
X_13458_ _06095_ _06145_ _06146_ vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__and3_1
XFILLER_51_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12409_ _05078_ _05080_ _05084_ _05101_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__or4_1
X_16177_ _07471_ _08787_ _08788_ _07697_ vssd1 vssd1 vccd1 vccd1 _08789_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_115_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13389_ _06042_ _06076_ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15128_ _07442_ vssd1 vssd1 vccd1 vccd1 _07742_ sky130_fd_sc_hd__buf_2
XFILLER_115_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15059_ _04936_ rbzero.wall_tracer.stepDistX\[0\] vssd1 vssd1 vccd1 vccd1 _07673_
+ sky130_fd_sc_hd__nand2_2
XFILLER_173_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19936_ _03116_ vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__clkinv_2
XFILLER_151_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19867_ _03109_ vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__clkinv_2
XFILLER_25_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18818_ _02520_ _02535_ _02536_ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__or3_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19798_ gpout0.vpos\[6\] _03096_ _03098_ _03031_ vssd1 vssd1 vccd1 vccd1 _01043_
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18749_ _02472_ rbzero.wall_tracer.rayAddendY\[3\] vssd1 vssd1 vccd1 vccd1 _02473_
+ sky130_fd_sc_hd__nand2_1
XFILLER_97_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20711_ net109 _00727_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.ss_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20642_ net66 _00658_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_189_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20573_ net101 _00589_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vinf sky130_fd_sc_hd__dfxtp_1
XFILLER_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21125_ _00174_ _01141_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21056_ _00105_ _01072_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20007_ _03123_ vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__clkinv_2
XFILLER_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _05346_ _05353_ _05448_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__mux2_1
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ rbzero.tex_g1\[46\] _04374_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__and2_1
XFILLER_243_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20909_ net61 _00925_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[46\] sky130_fd_sc_hd__dfxtp_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12691_ _05305_ _05256_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__nand2_1
XFILLER_226_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14430_ rbzero.wall_tracer.stepDistY\[-12\] _07118_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _07119_ sky130_fd_sc_hd__mux2_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _03957_ _04356_ _04357_ _04358_ _03920_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__o221a_1
XFILLER_230_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14361_ _07045_ _07049_ _05531_ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__mux2_1
XFILLER_168_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11573_ rbzero.debug_overlay.playerX\[-4\] _04242_ _04244_ rbzero.debug_overlay.playerX\[-1\]
+ _04290_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__a221o_1
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16100_ _08666_ _08682_ vssd1 vssd1 vccd1 vccd1 _08712_ sky130_fd_sc_hd__or2b_1
XFILLER_183_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 i_gpout2_sel[3] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_4
XFILLER_210_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13312_ _05958_ _06000_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__xor2_1
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17080_ _09460_ _09484_ _09620_ vssd1 vssd1 vccd1 vccd1 _09621_ sky130_fd_sc_hd__a21bo_1
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 i_gpout4_sel[2] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_4
X_10524_ _03445_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__clkbuf_4
X_14292_ _05593_ vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__buf_2
XFILLER_182_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16031_ _08473_ _08477_ vssd1 vssd1 vccd1 vccd1 _08644_ sky130_fd_sc_hd__and2_1
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13243_ _05904_ _05930_ _05931_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__o21a_1
XFILLER_202_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10455_ rbzero.tex_r1\[0\] rbzero.tex_r1\[1\] _03433_ vssd1 vssd1 vccd1 vccd1 _03441_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13174_ _05616_ _05728_ _05726_ _05611_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__o22a_1
XFILLER_48_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10386_ rbzero.tex_r1\[33\] rbzero.tex_r1\[34\] _03400_ vssd1 vssd1 vccd1 vccd1 _03405_
+ sky130_fd_sc_hd__mux2_1
XFILLER_184_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12125_ net32 net31 _04831_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__and3_1
XFILLER_124_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17982_ _01762_ _01763_ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__nand2_1
XFILLER_81_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19721_ rbzero.pov.ready_buffer\[41\] _03061_ _03063_ rbzero.debug_overlay.facingX\[-1\]
+ _03066_ vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__a221o_1
X_16933_ _08335_ _09200_ _07835_ vssd1 vssd1 vccd1 vccd1 _09475_ sky130_fd_sc_hd__o21ai_1
XFILLER_238_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12056_ net5 _04735_ _04760_ _04764_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a31o_1
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11007_ rbzero.map_rom.f3 vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__inv_2
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19652_ rbzero.debug_overlay.playerY\[-7\] _03016_ _03018_ _02978_ vssd1 vssd1 vccd1
+ vccd1 _00977_ sky130_fd_sc_hd__o211a_1
X_16864_ _08595_ _09166_ _09164_ _09405_ vssd1 vssd1 vccd1 vccd1 _09406_ sky130_fd_sc_hd__o31a_1
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18603_ _02335_ _05183_ _02326_ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__or3_1
X_15815_ _07616_ vssd1 vssd1 vccd1 vccd1 _08429_ sky130_fd_sc_hd__clkbuf_4
XFILLER_168_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16795_ _09339_ _09340_ vssd1 vssd1 vccd1 vccd1 _09341_ sky130_fd_sc_hd__and2b_1
X_19583_ _02956_ _02964_ _02965_ _02780_ vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__o211a_1
XFILLER_24_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15746_ _07468_ _08060_ vssd1 vssd1 vccd1 vccd1 _08360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18534_ _02247_ rbzero.wall_tracer.rayAddendX\[5\] vssd1 vssd1 vccd1 vccd1 _02278_
+ sky130_fd_sc_hd__or2_1
X_12958_ _05645_ _05634_ _05618_ _05646_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__a22oi_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11909_ _04611_ o_rgb[7] _04619_ net13 vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a211o_1
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15677_ _08251_ _08260_ vssd1 vssd1 vccd1 vccd1 _08291_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18465_ _02208_ _02213_ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__or2_1
X_12889_ _05314_ _05435_ _05430_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__mux2_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17416_ _09849_ _09855_ _09953_ vssd1 vssd1 vccd1 vccd1 _09954_ sky130_fd_sc_hd__a21oi_1
X_14628_ _07245_ _07280_ _07281_ _07251_ vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__o211a_1
X_18396_ _02148_ _02149_ _02147_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__nand3b_1
XFILLER_187_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17347_ _09759_ _09763_ _09757_ vssd1 vssd1 vccd1 vccd1 _09886_ sky130_fd_sc_hd__a21bo_1
XFILLER_109_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14559_ _07101_ _07228_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__nand2_2
XFILLER_187_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17278_ _09815_ _09816_ vssd1 vssd1 vccd1 vccd1 _09817_ sky130_fd_sc_hd__and2b_1
XFILLER_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16229_ _08822_ _08823_ vssd1 vssd1 vccd1 vccd1 _08840_ sky130_fd_sc_hd__or2_2
X_19017_ _02669_ vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19919_ _03115_ vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__clkinv_2
XFILLER_116_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20625_ net79 _00641_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20556_ net121 _00572_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20487_ net112 _00503_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10240_ rbzero.tex_b1\[38\] rbzero.tex_b1\[39\] _03322_ vssd1 vssd1 vccd1 vccd1 _03328_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21108_ _00157_ _01124_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_6868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout140 net141 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_2
XFILLER_134_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13930_ _06605_ _06617_ _06618_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__a21oi_1
XFILLER_43_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21039_ _00088_ _01055_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13861_ _06489_ _06549_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__and2_1
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15600_ _08191_ _08212_ _08213_ vssd1 vssd1 vccd1 vccd1 _08214_ sky130_fd_sc_hd__a21boi_2
XFILLER_210_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12812_ _05444_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__buf_2
XFILLER_41_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16580_ _08478_ _08928_ _07814_ vssd1 vssd1 vccd1 vccd1 _09189_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13792_ _06167_ _06173_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__nor2_1
XFILLER_76_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15531_ _08131_ _08144_ vssd1 vssd1 vccd1 vccd1 _08145_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12743_ _05431_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__buf_2
XFILLER_163_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18250_ _02021_ _02022_ _02023_ vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__o21ai_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15462_ _08021_ _08019_ _08020_ vssd1 vssd1 vccd1 vccd1 _08076_ sky130_fd_sc_hd__and3_1
X_12674_ _05362_ _05355_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__nand2_2
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _09615_ _09617_ vssd1 vssd1 vccd1 vccd1 _09741_ sky130_fd_sc_hd__or2b_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _07101_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__buf_4
XFILLER_141_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18181_ _01953_ _01960_ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11625_ _04340_ _04341_ _03942_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__mux2_1
XFILLER_204_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15393_ _07938_ _07939_ vssd1 vssd1 vccd1 vccd1 _08007_ sky130_fd_sc_hd__xnor2_2
XFILLER_180_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17132_ _09670_ _09671_ vssd1 vssd1 vccd1 vccd1 _09672_ sky130_fd_sc_hd__xor2_1
XFILLER_168_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14344_ _05432_ _06979_ _06983_ vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__and3_1
XFILLER_204_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11556_ _04269_ _04273_ gpout0.vpos\[5\] _04102_ _04246_ vssd1 vssd1 vccd1 vccd1
+ _04274_ sky130_fd_sc_hd__o2111a_1
XFILLER_102_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17063_ _07814_ _09462_ _09467_ _09603_ vssd1 vssd1 vccd1 vccd1 _09604_ sky130_fd_sc_hd__or4_1
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10507_ _03470_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__clkbuf_1
X_14275_ _06788_ _06963_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11487_ _03788_ _04202_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__nor2_1
X_16014_ _07814_ _07834_ vssd1 vssd1 vccd1 vccd1 _08627_ sky130_fd_sc_hd__nor2_1
X_13226_ _05913_ _05914_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10438_ rbzero.tex_r1\[8\] rbzero.tex_r1\[9\] _03422_ vssd1 vssd1 vccd1 vccd1 _03432_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_1262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13157_ _05747_ _05750_ _05751_ _05752_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__a22o_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ rbzero.tex_r1\[41\] rbzero.tex_r1\[42\] _03389_ vssd1 vssd1 vccd1 vccd1 _03396_
+ sky130_fd_sc_hd__mux2_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12108_ _04803_ _04815_ _04809_ _04779_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__o211a_1
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17965_ _01638_ _01639_ _09978_ _01637_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__o2bb2a_1
X_13088_ _05775_ _05776_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__and2_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19704_ _03057_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__clkbuf_2
X_16916_ _09202_ _09204_ _09456_ vssd1 vssd1 vccd1 vccd1 _09458_ sky130_fd_sc_hd__or3_1
XFILLER_239_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12039_ net3 _04718_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__and2b_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17896_ _01452_ _01455_ _01554_ vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__a21oi_1
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19635_ rbzero.debug_overlay.playerX\[5\] _03000_ _02835_ vssd1 vssd1 vccd1 vccd1
+ _03005_ sky130_fd_sc_hd__a21oi_1
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16847_ _09388_ vssd1 vssd1 vccd1 vccd1 _09389_ sky130_fd_sc_hd__buf_4
XFILLER_38_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19566_ rbzero.pov.sclk_buffer\[1\] rbzero.pov.sclk_buffer\[0\] _09243_ vssd1 vssd1
+ vccd1 vccd1 _02952_ sky130_fd_sc_hd__mux2_1
XFILLER_94_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16778_ rbzero.wall_tracer.trackDistX\[-6\] rbzero.wall_tracer.stepDistX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _09326_ sky130_fd_sc_hd__and2_1
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18517_ rbzero.debug_overlay.vplaneX\[0\] rbzero.debug_overlay.vplaneX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__and2_1
X_15729_ _08332_ _08342_ vssd1 vssd1 vccd1 vccd1 _08343_ sky130_fd_sc_hd__xnor2_1
XFILLER_248_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19497_ _02916_ vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18448_ rbzero.debug_overlay.vplaneX\[-5\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__or2_1
XFILLER_181_1258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18379_ _01916_ _02135_ _01996_ rbzero.wall_tracer.trackDistY\[10\] vssd1 vssd1 vccd1
+ vccd1 _00587_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_239_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20410_ net130 _00441_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_144_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21390_ net110 _01406_ vssd1 vssd1 vccd1 vccd1 gpout0.clk_div\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20341_ _02153_ _03271_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__xnor2_1
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20272_ _03125_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__buf_4
XFILLER_143_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11410_ rbzero.tex_r1\[61\] rbzero.tex_r1\[60\] _03935_ vssd1 vssd1 vccd1 vccd1 _04128_
+ sky130_fd_sc_hd__mux2_1
X_20608_ net90 _00624_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12390_ _05031_ _05032_ _05081_ _05082_ _05035_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__a221o_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11341_ _04055_ gpout0.hpos\[3\] gpout0.hpos\[2\] _04041_ _04059_ vssd1 vssd1 vccd1
+ vccd1 _04060_ sky130_fd_sc_hd__o221a_1
X_20539_ net139 _00555_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14060_ _06317_ _06634_ _06542_ _05767_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__o22a_1
XFILLER_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11272_ rbzero.tex_r0\[23\] rbzero.tex_r0\[22\] _03974_ vssd1 vssd1 vccd1 vccd1 _03991_
+ sky130_fd_sc_hd__mux2_1
XFILLER_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13011_ _05433_ _05606_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__nor2_2
XFILLER_238_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10223_ rbzero.tex_b1\[46\] rbzero.tex_b1\[47\] _03311_ vssd1 vssd1 vccd1 vccd1 _03319_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17750_ _09833_ _08531_ _08985_ _09571_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__o22a_1
X_14962_ _07567_ _07575_ vssd1 vssd1 vccd1 vccd1 _07576_ sky130_fd_sc_hd__or2_1
XFILLER_43_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16701_ rbzero.traced_texa\[3\] _09264_ _09265_ rbzero.wall_tracer.visualWallDist\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__a22o_1
XFILLER_59_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13913_ _06583_ _06601_ vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__xnor2_1
XFILLER_235_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17681_ _08241_ _09463_ _09962_ _01465_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__o31a_1
X_14893_ _04928_ rbzero.wall_tracer.stepDistX\[-9\] _07505_ _07506_ vssd1 vssd1 vccd1
+ vccd1 _07507_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_207_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19420_ rbzero.pov.spi_buffer\[8\] rbzero.pov.spi_buffer\[9\] _02866_ vssd1 vssd1
+ vccd1 vccd1 _02876_ sky130_fd_sc_hd__mux2_1
X_13844_ _06524_ _06525_ _06531_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__a21oi_1
X_16632_ _09108_ _09240_ vssd1 vssd1 vccd1 vccd1 _09241_ sky130_fd_sc_hd__xnor2_1
XFILLER_207_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19351_ _02858_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__clkinv_2
X_16563_ _07890_ _07834_ vssd1 vssd1 vccd1 vccd1 _09172_ sky130_fd_sc_hd__nor2_1
X_13775_ _06115_ _06320_ _06461_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__a21o_1
XFILLER_188_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10987_ rbzero.tex_b0\[6\] rbzero.tex_b0\[5\] _03715_ vssd1 vssd1 vccd1 vccd1 _03722_
+ sky130_fd_sc_hd__mux2_1
XFILLER_203_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18302_ _04953_ _02001_ _02069_ vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__a21oi_1
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15514_ _08048_ _08127_ vssd1 vssd1 vccd1 vccd1 _08128_ sky130_fd_sc_hd__xor2_1
X_12726_ _05348_ _05411_ _05414_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__and3b_1
X_16494_ _08585_ _09103_ vssd1 vssd1 vccd1 vccd1 _09104_ sky130_fd_sc_hd__xnor2_1
X_19282_ rbzero.spi_registers.new_vshift\[0\] rbzero.spi_registers.spi_buffer\[0\]
+ _02825_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__mux2_1
XFILLER_188_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15445_ _04936_ rbzero.wall_tracer.stepDistX\[-12\] _07633_ vssd1 vssd1 vccd1 vccd1
+ _08059_ sky130_fd_sc_hd__a21boi_4
X_18233_ rbzero.wall_tracer.trackDistY\[-10\] rbzero.wall_tracer.stepDistY\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__and2_1
XFILLER_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12657_ _05340_ _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__xor2_4
XFILLER_19_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11608_ rbzero.tex_g0\[6\] _04013_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__and2_1
X_18164_ _01942_ _01943_ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__xor2_1
X_15376_ _07567_ _07986_ _07989_ _07987_ vssd1 vssd1 vccd1 vccd1 _07990_ sky130_fd_sc_hd__o31a_1
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12588_ _05199_ _05204_ _05271_ _05276_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__or4_2
XFILLER_89_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17115_ _09654_ vssd1 vssd1 vccd1 vccd1 _09655_ sky130_fd_sc_hd__inv_2
X_14327_ _07011_ _07015_ vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__or2_1
XFILLER_15_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18095_ _01874_ _01875_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11539_ rbzero.debug_overlay.vplaneX\[-7\] _04238_ _04254_ _04256_ vssd1 vssd1 vccd1
+ vccd1 _04257_ sky130_fd_sc_hd__a211o_1
XFILLER_89_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17046_ _09569_ _09585_ vssd1 vssd1 vccd1 vccd1 _09587_ sky130_fd_sc_hd__or2_1
XFILLER_183_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14258_ _06934_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__inv_2
XFILLER_99_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13209_ _05894_ _05897_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__or2b_1
XFILLER_171_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14189_ _06835_ _06837_ _06809_ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__a21oi_1
XFILLER_174_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18997_ rbzero.pov.spi_buffer\[46\] rbzero.pov.ready_buffer\[46\] _02651_ vssd1 vssd1
+ vccd1 vccd1 _02659_ sky130_fd_sc_hd__mux2_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _09861_ _09989_ _01621_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__nor3_2
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17879_ _10056_ _08724_ _01534_ _01536_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__o31a_1
XFILLER_96_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19618_ rbzero.debug_overlay.playerX\[2\] rbzero.debug_overlay.playerX\[1\] _02982_
+ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__or3_1
XFILLER_54_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20890_ net66 _00906_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_241_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19549_ _02943_ vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__clkbuf_1
XFILLER_228_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21373_ _00396_ _01389_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20324_ gpout0.clk_div\[0\] gpout0.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__nand2_1
XFILLER_135_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20255_ _03254_ vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__clkinv_2
XFILLER_153_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20186_ _03209_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__inv_2
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10910_ _03681_ vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__clkbuf_1
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ rbzero.row_render.texu\[0\] _03289_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__or2b_1
XFILLER_217_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10841_ _03645_ vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13560_ _06247_ _06248_ vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__nand2_1
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10772_ _03609_ vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ _03816_ _05080_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__nand2_1
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13491_ _05856_ _05870_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__and2b_1
XFILLER_164_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15230_ _07840_ _07843_ vssd1 vssd1 vccd1 vccd1 _07844_ sky130_fd_sc_hd__nor2_1
XFILLER_185_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12442_ _05131_ _05132_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__nand2_1
XFILLER_90_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15161_ _07767_ _07769_ _07766_ vssd1 vssd1 vccd1 vccd1 _07775_ sky130_fd_sc_hd__a21o_1
XFILLER_176_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12373_ rbzero.wall_tracer.rayAddendY\[10\] rbzero.wall_tracer.rayAddendY\[9\] rbzero.debug_overlay.facingY\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__o21ai_1
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14112_ _06435_ _06483_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__nor2_1
XFILLER_165_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11324_ _04041_ _04042_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__nand2_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15092_ _07342_ _05100_ _07705_ _07346_ vssd1 vssd1 vccd1 vccd1 _07706_ sky130_fd_sc_hd__o211a_1
XFILLER_153_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14043_ _06707_ _06731_ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__xor2_2
X_18920_ rbzero.pov.spi_buffer\[9\] rbzero.pov.ready_buffer\[9\] _02618_ vssd1 vssd1
+ vccd1 vccd1 _02619_ sky130_fd_sc_hd__mux2_1
XTAP_7130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11255_ _03903_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__buf_4
XTAP_7141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10206_ rbzero.tex_b1\[54\] rbzero.tex_b1\[55\] _03300_ vssd1 vssd1 vccd1 vccd1 _03310_
+ sky130_fd_sc_hd__mux2_1
XFILLER_175_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18851_ _02510_ _03818_ _02567_ vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__or3_1
XTAP_6440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11186_ rbzero.tex_r0\[49\] rbzero.tex_r0\[48\] _03904_ vssd1 vssd1 vccd1 vccd1 _03905_
+ sky130_fd_sc_hd__mux2_1
XTAP_6451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17802_ _01472_ _01473_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__nand2_1
XFILLER_67_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18782_ _02502_ _02503_ vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__xnor2_1
XTAP_6495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15994_ _08605_ _08606_ vssd1 vssd1 vccd1 vccd1 _08607_ sky130_fd_sc_hd__xnor2_1
XTAP_5750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17733_ _08750_ _09115_ _10165_ _10166_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__o31a_1
XTAP_5783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14945_ _07558_ rbzero.debug_overlay.playerY\[-1\] _05114_ vssd1 vssd1 vccd1 vccd1
+ _07559_ sky130_fd_sc_hd__mux2_1
XTAP_5794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17664_ _10103_ _10105_ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__nor2_1
XFILLER_208_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14876_ _07488_ _07489_ vssd1 vssd1 vccd1 vccd1 _07490_ sky130_fd_sc_hd__nand2_1
XFILLER_211_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19403_ _02867_ vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__clkbuf_1
XFILLER_223_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16615_ _09081_ _09083_ vssd1 vssd1 vccd1 vccd1 _09224_ sky130_fd_sc_hd__and2_1
XFILLER_169_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13827_ _06515_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__clkbuf_2
X_17595_ _10130_ _10131_ vssd1 vssd1 vccd1 vccd1 _10132_ sky130_fd_sc_hd__xor2_1
XFILLER_189_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19334_ _02856_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__clkinv_2
X_16546_ _09140_ _09154_ vssd1 vssd1 vccd1 vccd1 _09155_ sky130_fd_sc_hd__xnor2_1
X_13758_ _06432_ _06445_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__and2_1
XFILLER_245_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12709_ _05361_ _05351_ _05335_ _05344_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__or4_1
XFILLER_143_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19265_ rbzero.spi_registers.new_other\[3\] rbzero.spi_registers.spi_buffer\[3\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__mux2_1
XFILLER_231_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16477_ _09083_ _09084_ _09086_ vssd1 vssd1 vccd1 vccd1 _09087_ sky130_fd_sc_hd__nand3_1
XFILLER_182_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13689_ _06230_ _06321_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__and2_1
XFILLER_206_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18216_ _03797_ _08629_ _05027_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__o21a_4
XFILLER_176_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15428_ _08037_ _08040_ _08041_ vssd1 vssd1 vccd1 vccd1 _08042_ sky130_fd_sc_hd__a21boi_1
XFILLER_31_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19196_ rbzero.spi_registers.vshift\[1\] _02774_ _02777_ _02738_ vssd1 vssd1 vccd1
+ vccd1 _00762_ sky130_fd_sc_hd__o211a_1
XFILLER_191_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18147_ _01925_ _01926_ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__xnor2_1
X_15359_ _07969_ _07972_ vssd1 vssd1 vccd1 vccd1 _07973_ sky130_fd_sc_hd__xnor2_2
XFILLER_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18078_ _01857_ _01858_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__or2b_1
XFILLER_160_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17029_ _07591_ _07790_ _07672_ _07817_ vssd1 vssd1 vccd1 vccd1 _09570_ sky130_fd_sc_hd__or4_1
XFILLER_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20040_ _03127_ vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__clkinv_2
XFILLER_193_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20942_ net85 _00958_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_226_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20873_ net56 _00889_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21356_ _00379_ _01372_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20307_ _02855_ vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__clkinv_2
XFILLER_190_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21287_ _00336_ _01303_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[63\] sky130_fd_sc_hd__dfxtp_1
X_11040_ rbzero.otherx\[1\] _03735_ rbzero.map_rom.i_row\[4\] _03766_ _03767_ vssd1
+ vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__o221a_1
XFILLER_89_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20238_ _03251_ _03252_ rbzero.texV\[11\] _03003_ vssd1 vssd1 vccd1 vccd1 _01329_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20169_ _03189_ _03191_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__nand2_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _05604_ _05622_ _05679_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__or3b_1
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14730_ _07339_ _07340_ _07343_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__mux2_1
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11942_ net14 net13 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__nor2_1
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14661_ rbzero.wall_tracer.trackDistX\[10\] rbzero.wall_tracer.trackDistY\[10\] _05025_
+ vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__mux2_1
XFILLER_189_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _03896_ _04535_ _04553_ _04569_ _04586_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__o32a_1
XFILLER_73_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16400_ _08976_ _08977_ _09009_ vssd1 vssd1 vccd1 vccd1 _09010_ sky130_fd_sc_hd__a21o_1
XFILLER_207_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13612_ _06214_ _06254_ _06256_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__a21o_1
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10824_ _03636_ vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17380_ _08507_ _09114_ vssd1 vssd1 vccd1 vccd1 _09918_ sky130_fd_sc_hd__nor2_1
X_14592_ _04968_ _07246_ _07253_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__o21ai_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16331_ _08802_ _08804_ vssd1 vssd1 vccd1 vccd1 _08942_ sky130_fd_sc_hd__nor2_1
X_13543_ _05624_ _05610_ _05749_ vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__o21ai_1
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10755_ rbzero.tex_g0\[52\] rbzero.tex_g0\[51\] _03593_ vssd1 vssd1 vccd1 vccd1 _03600_
+ sky130_fd_sc_hd__mux2_1
XFILLER_198_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16262_ _08729_ _08738_ _08872_ vssd1 vssd1 vccd1 vccd1 _08873_ sky130_fd_sc_hd__a21oi_1
XFILLER_158_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19050_ _02686_ vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13474_ _05881_ _06162_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__xnor2_1
X_10686_ _03564_ vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18001_ _07618_ _07827_ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__nor2_1
XFILLER_199_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15213_ _07824_ vssd1 vssd1 vccd1 vccd1 _07827_ sky130_fd_sc_hd__clkbuf_4
XFILLER_185_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12425_ _03743_ _05117_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__xnor2_1
X_16193_ _08802_ _08804_ vssd1 vssd1 vccd1 vccd1 _08805_ sky130_fd_sc_hd__xor2_1
XFILLER_200_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15144_ _07720_ _07721_ vssd1 vssd1 vccd1 vccd1 _07758_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12356_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__nand2_1
XFILLER_5_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ _03879_ _03894_ _03895_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__nor3_4
XFILLER_99_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15075_ _07101_ _07216_ vssd1 vssd1 vccd1 vccd1 _07689_ sky130_fd_sc_hd__and2_1
XFILLER_142_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19952_ _03118_ vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__clkinv_2
X_12287_ _04980_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__inv_2
XFILLER_141_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14026_ _06407_ _06691_ _06692_ vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__a21bo_1
XFILLER_113_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18903_ rbzero.pov.spi_buffer\[1\] rbzero.pov.ready_buffer\[1\] _02608_ vssd1 vssd1
+ vccd1 vccd1 _02610_ sky130_fd_sc_hd__mux2_1
X_11238_ _03909_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__buf_4
XFILLER_136_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19883_ _03111_ vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__clkinv_2
XFILLER_218_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18834_ _03818_ _02551_ _02552_ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__or3_1
XTAP_6270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11169_ rbzero.traced_texVinit\[9\] rbzero.texV\[9\] _03880_ _03881_ _03887_ vssd1
+ vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__a41o_1
XTAP_6281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18765_ _02473_ _02478_ _02487_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__a21oi_1
X_15977_ _08512_ _08520_ _08519_ vssd1 vssd1 vccd1 vccd1 _08590_ sky130_fd_sc_hd__a21o_1
XTAP_5580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17716_ _10020_ _10145_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__nor2_1
XFILLER_208_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14928_ _07356_ _07536_ _07541_ vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__o21ai_4
XFILLER_3_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18696_ _02422_ _02423_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__nand2_1
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17647_ _07619_ _07663_ _08536_ _07651_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_224_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14859_ _07470_ _07442_ _07471_ _07472_ vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__o22ai_1
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17578_ _09182_ _09603_ _10112_ _10113_ vssd1 vssd1 vccd1 vccd1 _10115_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_223_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19317_ rbzero.pov.spi_counter\[4\] rbzero.pov.spi_counter\[3\] _02846_ vssd1 vssd1
+ vccd1 vccd1 _02849_ sky130_fd_sc_hd__and3_1
X_16529_ _09128_ _09137_ vssd1 vssd1 vccd1 vccd1 _09138_ sky130_fd_sc_hd__nand2_1
XFILLER_189_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19248_ _02807_ vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19179_ rbzero.color_floor\[1\] _02763_ _02766_ vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__a21o_1
XFILLER_247_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21210_ _00259_ _01226_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21141_ _00190_ _01157_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21072_ _00121_ _01088_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_232_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20023_ _03124_ vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__clkinv_2
XFILLER_86_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20925_ net75 _00941_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[62\] sky130_fd_sc_hd__dfxtp_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20856_ _00074_ _00872_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_230_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20787_ net102 _00803_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10540_ _03487_ vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10471_ _03451_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12210_ net37 _04910_ _04915_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__and3b_1
XFILLER_202_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13190_ _05839_ _05878_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__xor2_1
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12141_ _04840_ net27 vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__and2_1
XFILLER_159_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21339_ _00362_ _01355_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12072_ net22 net23 net24 vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__a21o_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15900_ _07742_ _07890_ _07800_ _07469_ vssd1 vssd1 vccd1 vccd1 _08514_ sky130_fd_sc_hd__o22ai_1
X_11023_ _03736_ rbzero.map_rom.f1 rbzero.map_rom.i_col\[4\] vssd1 vssd1 vccd1 vccd1
+ _03751_ sky130_fd_sc_hd__and3_1
XFILLER_133_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16880_ _09420_ _09421_ vssd1 vssd1 vccd1 vccd1 _09422_ sky130_fd_sc_hd__nand2_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15831_ _08411_ _08441_ _08355_ _08442_ _08444_ vssd1 vssd1 vccd1 vccd1 _08445_ sky130_fd_sc_hd__o2111a_1
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ _02274_ rbzero.debug_overlay.vplaneX\[-3\] _02291_ _02292_ vssd1 vssd1 vccd1
+ vccd1 _02293_ sky130_fd_sc_hd__o22ai_1
XFILLER_218_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15762_ _08360_ _08362_ _08361_ vssd1 vssd1 vccd1 vccd1 _08376_ sky130_fd_sc_hd__a21boi_1
X_12974_ _05662_ _05658_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__or2b_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ _09779_ _09781_ _09911_ _09909_ vssd1 vssd1 vccd1 vccd1 _10038_ sky130_fd_sc_hd__a31o_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ rbzero.wall_tracer.stepDistX\[11\] _07243_ _04931_ vssd1 vssd1 vccd1 vccd1
+ _07331_ sky130_fd_sc_hd__mux2_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11925_ net12 _04635_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__or2_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18481_ _02210_ _02228_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__xnor2_1
XFILLER_233_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15693_ _08291_ _08305_ vssd1 vssd1 vccd1 vccd1 _08307_ sky130_fd_sc_hd__or2b_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _09967_ _09969_ vssd1 vssd1 vccd1 vccd1 _09970_ sky130_fd_sc_hd__xor2_1
XFILLER_2_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14644_ rbzero.wall_tracer.visualWallDist\[4\] _07253_ _07290_ _07292_ _07266_ vssd1
+ vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__o221a_1
X_11856_ rbzero.tex_b1\[15\] rbzero.tex_b1\[14\] _04544_ vssd1 vssd1 vccd1 vccd1 _04570_
+ sky130_fd_sc_hd__mux2_1
XFILLER_205_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10807_ rbzero.tex_g0\[28\] rbzero.tex_g0\[27\] _03627_ vssd1 vssd1 vccd1 vccd1 _03628_
+ sky130_fd_sc_hd__mux2_1
X_17363_ _09791_ _09823_ vssd1 vssd1 vccd1 vccd1 _09901_ sky130_fd_sc_hd__nand2_1
X_14575_ rbzero.wall_tracer.stepDistY\[10\] _07241_ _04925_ vssd1 vssd1 vccd1 vccd1
+ _07242_ sky130_fd_sc_hd__mux2_1
XFILLER_183_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11787_ rbzero.tex_b0\[5\] rbzero.tex_b0\[4\] _04001_ vssd1 vssd1 vccd1 vccd1 _04502_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19102_ rbzero.spi_registers.sclk_buffer\[2\] rbzero.spi_registers.sclk_buffer\[1\]
+ _09243_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__mux2_1
XFILLER_92_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16314_ _07826_ _08917_ _08923_ _07471_ vssd1 vssd1 vccd1 vccd1 _08925_ sky130_fd_sc_hd__o22a_1
XFILLER_186_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13526_ _05872_ _06179_ _06213_ vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__and3_1
X_10738_ rbzero.tex_g0\[60\] rbzero.tex_g0\[59\] _03512_ vssd1 vssd1 vccd1 vccd1 _03591_
+ sky130_fd_sc_hd__mux2_1
X_17294_ _07472_ vssd1 vssd1 vccd1 vccd1 _09833_ sky130_fd_sc_hd__buf_2
XFILLER_158_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19033_ rbzero.pov.spi_buffer\[63\] rbzero.pov.ready_buffer\[63\] _02673_ vssd1 vssd1
+ vccd1 vccd1 _02678_ sky130_fd_sc_hd__mux2_1
X_16245_ _07878_ _08718_ _08855_ _07521_ vssd1 vssd1 vccd1 vccd1 _08856_ sky130_fd_sc_hd__a2bb2o_1
X_13457_ _06093_ _06089_ _06092_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__nand3_1
XFILLER_220_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10669_ _03555_ vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__clkbuf_1
X_12408_ _05085_ _05089_ _05098_ _05100_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__or4_1
X_16176_ _07696_ _08640_ vssd1 vssd1 vccd1 vccd1 _08788_ sky130_fd_sc_hd__nand2_2
XFILLER_220_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13388_ _05625_ _05660_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__or2_1
XFILLER_217_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15127_ _07715_ _07740_ vssd1 vssd1 vccd1 vccd1 _07741_ sky130_fd_sc_hd__xor2_1
X_12339_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__or2_1
XFILLER_47_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15058_ _03794_ _07670_ _07671_ _07356_ vssd1 vssd1 vccd1 vccd1 _07672_ sky130_fd_sc_hd__a211o_2
X_19935_ _03116_ vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__clkinv_2
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14009_ _06310_ _06483_ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__nor2_1
XFILLER_123_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19866_ _03109_ vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__clkinv_2
XFILLER_60_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18817_ _02535_ _02536_ _02520_ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__o21ai_1
XFILLER_233_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19797_ gpout0.vpos\[6\] _03096_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__nand2_1
XFILLER_37_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18748_ rbzero.debug_overlay.vplaneY\[10\] vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__buf_2
XFILLER_243_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18679_ _04260_ rbzero.wall_tracer.rayAddendY\[-2\] vssd1 vssd1 vccd1 vccd1 _02408_
+ sky130_fd_sc_hd__nand2_1
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20710_ net85 _00726_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.mosi sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20641_ net56 _00657_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_189_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20572_ net124 _00588_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21124_ _00173_ _01140_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21055_ _00104_ _01071_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20006_ _03123_ vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__clkinv_2
XFILLER_219_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11710_ rbzero.tex_g1\[45\] rbzero.tex_g1\[44\] _03962_ vssd1 vssd1 vccd1 vccd1 _04426_
+ sky130_fd_sc_hd__mux2_1
XFILLER_226_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20908_ net61 _00924_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[45\] sky130_fd_sc_hd__dfxtp_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _05378_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__inv_2
XFILLER_128_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11641_ rbzero.tex_g0\[47\] _04142_ _04144_ _03915_ vssd1 vssd1 vccd1 vccd1 _04358_
+ sky130_fd_sc_hd__a31o_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20839_ _00057_ _00855_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14360_ _06987_ _07048_ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__nor2_1
XFILLER_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11572_ rbzero.debug_overlay.playerX\[2\] _04235_ _04278_ rbzero.debug_overlay.playerX\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__a22o_1
XFILLER_122_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13311_ _05914_ _05957_ _05960_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__o21ba_1
XFILLER_122_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput19 i_gpout2_sel[4] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_6
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10523_ _03478_ vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14291_ _06368_ _06979_ vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__xor2_2
XFILLER_13_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16030_ _08641_ _08642_ vssd1 vssd1 vccd1 vccd1 _08643_ sky130_fd_sc_hd__xnor2_1
XFILLER_196_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13242_ _05905_ _05929_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__or2_1
XFILLER_196_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10454_ _03440_ vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13173_ _05607_ _05861_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__or2_1
XFILLER_170_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10385_ _03404_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_237_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12124_ net28 net29 net30 vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a21o_1
XFILLER_124_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17981_ _09429_ _09373_ _01761_ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__o21ai_1
XFILLER_111_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19720_ rbzero.pov.ready_buffer\[40\] _03061_ _03063_ rbzero.debug_overlay.facingX\[-2\]
+ _03066_ vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__a221o_1
X_16932_ _07835_ _08335_ _09200_ vssd1 vssd1 vccd1 vccd1 _09474_ sky130_fd_sc_hd__or3_1
X_12055_ _04719_ _04762_ _04763_ _04743_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__a22o_1
XFILLER_172_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11006_ _03733_ rbzero.map_rom.a6 vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__nand2_1
X_19651_ rbzero.pov.ready_buffer\[46\] _02836_ _03008_ _03017_ vssd1 vssd1 vccd1 vccd1
+ _03018_ sky130_fd_sc_hd__a211o_1
X_16863_ _08067_ _07685_ _09028_ vssd1 vssd1 vccd1 vccd1 _09405_ sky130_fd_sc_hd__or3b_1
XFILLER_120_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18602_ rbzero.wall_tracer.rayAddendX\[10\] _02158_ _02336_ _02340_ vssd1 vssd1 vccd1
+ vccd1 _00605_ sky130_fd_sc_hd__a211o_1
XFILLER_19_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15814_ _07878_ _08398_ _08425_ vssd1 vssd1 vccd1 vccd1 _08428_ sky130_fd_sc_hd__o21a_1
XFILLER_237_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19582_ _07431_ _02960_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__nand2_1
XFILLER_24_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16794_ rbzero.wall_tracer.trackDistX\[-4\] rbzero.wall_tracer.stepDistX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _09340_ sky130_fd_sc_hd__nand2_1
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18533_ _02247_ rbzero.wall_tracer.rayAddendX\[5\] vssd1 vssd1 vccd1 vccd1 _02277_
+ sky130_fd_sc_hd__nand2_1
X_15745_ _08341_ _08339_ _08340_ vssd1 vssd1 vccd1 vccd1 _08359_ sky130_fd_sc_hd__a21o_1
XFILLER_52_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12957_ _05611_ _05616_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__nand2_1
XFILLER_92_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18464_ _02211_ _02212_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__and2_1
X_11908_ _04611_ _04118_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__nor2_1
XFILLER_206_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15676_ _08280_ _08289_ vssd1 vssd1 vccd1 vccd1 _08290_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _05481_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__buf_2
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _09850_ _09854_ vssd1 vssd1 vccd1 vccd1 _09953_ sky130_fd_sc_hd__nor2_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14627_ rbzero.wall_tracer.visualWallDist\[-1\] _07252_ vssd1 vssd1 vccd1 vccd1 _07281_
+ sky130_fd_sc_hd__or2_1
XFILLER_21_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11839_ _03949_ _04539_ _04543_ _04552_ _03984_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__o311a_1
X_18395_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.wall_tracer.rayAddendX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__or2_1
XFILLER_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17346_ _09883_ _09884_ vssd1 vssd1 vccd1 vccd1 _09885_ sky130_fd_sc_hd__or2b_2
XFILLER_193_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14558_ _07007_ _07078_ _07214_ _07227_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__a22o_1
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13509_ _05692_ _05722_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__nand2_1
XFILLER_105_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17277_ _09809_ _09814_ vssd1 vssd1 vccd1 vccd1 _09816_ sky130_fd_sc_hd__nand2_1
XFILLER_186_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14489_ rbzero.wall_tracer.stepDistY\[-7\] _07172_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _07173_ sky130_fd_sc_hd__mux2_1
XFILLER_220_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19016_ rbzero.pov.spi_buffer\[55\] rbzero.pov.ready_buffer\[55\] _02662_ vssd1 vssd1
+ vccd1 vccd1 _02669_ sky130_fd_sc_hd__mux2_1
X_16228_ _08710_ _08827_ _08825_ vssd1 vssd1 vccd1 vccd1 _08839_ sky130_fd_sc_hd__a21bo_1
XFILLER_179_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16159_ _07964_ vssd1 vssd1 vccd1 vccd1 _08771_ sky130_fd_sc_hd__clkbuf_4
XFILLER_154_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19918_ _03115_ vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__clkinv_2
XFILLER_111_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19849_ _03108_ vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__clkinv_2
XFILLER_69_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20624_ net54 _00640_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20555_ net120 _00571_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20486_ net112 _00502_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21107_ _00156_ _01123_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout130 net140 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_2
XTAP_6869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout141 net1 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_4
XFILLER_134_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21038_ _00087_ _01054_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13860_ _06478_ _06488_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__nand2_1
XFILLER_210_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12811_ _05493_ _05498_ _05499_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__mux2_1
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13791_ _06479_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__inv_2
XFILLER_74_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15530_ _08133_ _08142_ _08143_ vssd1 vssd1 vccd1 vccd1 _08144_ sky130_fd_sc_hd__a21o_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _05430_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__buf_2
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15461_ _08023_ _08024_ vssd1 vssd1 vccd1 vccd1 _08075_ sky130_fd_sc_hd__xnor2_1
X_12673_ _05350_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__inv_2
XFILLER_163_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17200_ _09727_ _09739_ vssd1 vssd1 vccd1 vccd1 _09740_ sky130_fd_sc_hd__xnor2_1
XFILLER_230_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14412_ _07100_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__clkbuf_4
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11624_ rbzero.tex_g0\[53\] rbzero.tex_g0\[52\] _03935_ vssd1 vssd1 vccd1 vccd1 _04341_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18180_ _01956_ _01959_ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__xnor2_1
XFILLER_175_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15392_ _07942_ _07943_ _07944_ _07474_ vssd1 vssd1 vccd1 vccd1 _08006_ sky130_fd_sc_hd__a22o_1
XFILLER_169_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17131_ _08596_ _08724_ vssd1 vssd1 vccd1 vccd1 _09671_ sky130_fd_sc_hd__nor2_1
XFILLER_15_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14343_ _06981_ _06992_ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__and2_1
XFILLER_141_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11555_ rbzero.debug_overlay.facingY\[10\] _04236_ _04272_ vssd1 vssd1 vccd1 vccd1
+ _04273_ sky130_fd_sc_hd__a21o_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10506_ rbzero.tex_r0\[43\] rbzero.tex_r0\[42\] _03468_ vssd1 vssd1 vccd1 vccd1 _03470_
+ sky130_fd_sc_hd__mux2_1
XFILLER_221_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17062_ _09602_ vssd1 vssd1 vccd1 vccd1 _09603_ sky130_fd_sc_hd__clkbuf_4
X_14274_ _06782_ _06841_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__nor2_1
XFILLER_183_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11486_ _03788_ _04202_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__nand2_1
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16013_ _08624_ _08625_ vssd1 vssd1 vccd1 vccd1 _08626_ sky130_fd_sc_hd__and2_1
X_13225_ _05591_ _05627_ _05657_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__or3_1
X_10437_ _03431_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13156_ _05401_ _05738_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__nand2_1
XFILLER_174_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _03395_ vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ net46 _04798_ _04799_ _04702_ _04814_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__a221o_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ _01744_ _01745_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__xor2_1
X_13087_ _05769_ _05770_ _05774_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__or3_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ rbzero.tex_b1\[10\] rbzero.tex_b1\[11\] _03355_ vssd1 vssd1 vccd1 vccd1 _03359_
+ sky130_fd_sc_hd__mux2_1
XFILLER_239_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19703_ rbzero.pov.ready _02720_ _02833_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__and3_1
XFILLER_78_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16915_ _09202_ _09204_ _09456_ vssd1 vssd1 vccd1 vccd1 _09457_ sky130_fd_sc_hd__o21ai_1
X_12038_ _04718_ _03292_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__nor2_1
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17895_ _01669_ _01677_ vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19634_ rbzero.debug_overlay.playerX\[5\] _03001_ vssd1 vssd1 vccd1 vccd1 _03004_
+ sky130_fd_sc_hd__or2_1
X_16846_ rbzero.wall_tracer.visualWallDist\[11\] _03796_ _04929_ vssd1 vssd1 vccd1
+ vccd1 _09388_ sky130_fd_sc_hd__and3_1
XFILLER_4_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19565_ _02951_ vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__clkbuf_1
X_16777_ rbzero.wall_tracer.trackDistX\[-6\] rbzero.wall_tracer.stepDistX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _09325_ sky130_fd_sc_hd__nor2_1
XFILLER_4_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13989_ _06659_ _06677_ vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__xor2_1
XFILLER_209_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18516_ rbzero.debug_overlay.vplaneX\[0\] rbzero.debug_overlay.vplaneX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__nor2_1
XFILLER_206_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15728_ _08339_ _08340_ _08341_ vssd1 vssd1 vccd1 vccd1 _08342_ sky130_fd_sc_hd__a21bo_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19496_ rbzero.pov.spi_buffer\[44\] rbzero.pov.spi_buffer\[45\] _02910_ vssd1 vssd1
+ vccd1 vccd1 _02916_ sky130_fd_sc_hd__mux2_1
XFILLER_206_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18447_ _03810_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__clkbuf_4
X_15659_ _07467_ _07593_ vssd1 vssd1 vccd1 vccd1 _08273_ sky130_fd_sc_hd__or2_1
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18378_ _02133_ _02134_ _02039_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__o21a_1
XFILLER_193_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17329_ _09727_ _09739_ _09867_ vssd1 vssd1 vccd1 vccd1 _09868_ sky130_fd_sc_hd__a21o_1
XFILLER_147_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20340_ rbzero.debug_overlay.vplaneX\[-6\] rbzero.wall_tracer.rayAddendX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20271_ _03255_ vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__clkinv_2
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20607_ net90 _00623_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11340_ _04041_ gpout0.hpos\[2\] gpout0.hpos\[1\] _04056_ _04058_ vssd1 vssd1 vccd1
+ vccd1 _04059_ sky130_fd_sc_hd__a221o_1
X_20538_ net135 _00554_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11271_ rbzero.tex_r0\[21\] rbzero.tex_r0\[20\] _03974_ vssd1 vssd1 vccd1 vccd1 _03990_
+ sky130_fd_sc_hd__mux2_1
XFILLER_106_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20469_ net119 _00485_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ _05671_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__clkinv_2
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10222_ _03318_ vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14961_ _07574_ vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__buf_2
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16700_ rbzero.traced_texa\[2\] _09264_ _09265_ rbzero.wall_tracer.visualWallDist\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__a22o_1
XFILLER_248_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13912_ _06585_ _06600_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__xor2_1
XFILLER_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17680_ _10101_ _10102_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__nand2_1
XTAP_5987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14892_ _07408_ rbzero.wall_tracer.stepDistY\[-9\] _07352_ vssd1 vssd1 vccd1 vccd1
+ _07506_ sky130_fd_sc_hd__a21oi_1
XFILLER_169_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16631_ _09237_ _09239_ vssd1 vssd1 vccd1 vccd1 _09240_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13843_ _06524_ _06525_ _06531_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__and3_1
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19350_ _02858_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__clkinv_2
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16562_ _07751_ _08636_ vssd1 vssd1 vccd1 vccd1 _09171_ sky130_fd_sc_hd__and2b_1
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13774_ _06266_ _06343_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__nor2_1
X_10986_ _03721_ vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18301_ _09345_ _02067_ _02068_ _09361_ _01995_ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__o311a_1
XFILLER_71_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15513_ _08045_ _08047_ _08049_ vssd1 vssd1 vccd1 vccd1 _08127_ sky130_fd_sc_hd__o21ba_1
XFILLER_128_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12725_ _05391_ _05314_ _05318_ _05413_ _05307_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__o311a_1
XFILLER_43_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19281_ _03442_ _02824_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__nor2_4
XFILLER_231_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16493_ _09101_ _09102_ vssd1 vssd1 vccd1 vccd1 _09103_ sky130_fd_sc_hd__nand2_1
XFILLER_231_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18232_ rbzero.wall_tracer.trackDistY\[-10\] rbzero.wall_tracer.stepDistY\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__nor2_1
X_15444_ _08057_ _07989_ vssd1 vssd1 vccd1 vccd1 _08058_ sky130_fd_sc_hd__xor2_1
XFILLER_188_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12656_ _05338_ _05339_ _05341_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__a21o_1
XFILLER_175_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18163_ _08735_ _08645_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__nor2_1
X_11607_ rbzero.tex_g0\[5\] rbzero.tex_g0\[4\] _03936_ vssd1 vssd1 vccd1 vccd1 _04324_
+ sky130_fd_sc_hd__mux2_1
X_15375_ _07987_ _07988_ vssd1 vssd1 vccd1 vccd1 _07989_ sky130_fd_sc_hd__nand2_1
X_12587_ _03789_ _05273_ _05275_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__a21bo_2
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17114_ _08510_ _08852_ _09529_ _09533_ vssd1 vssd1 vccd1 vccd1 _09654_ sky130_fd_sc_hd__o31a_1
XFILLER_89_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14326_ _05431_ _07014_ vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__and2_1
XFILLER_144_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18094_ _08645_ _08671_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__nor2_1
XFILLER_141_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11538_ rbzero.debug_overlay.vplaneX\[-8\] _04218_ _04244_ rbzero.debug_overlay.vplaneX\[-1\]
+ _04255_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__a221o_1
XFILLER_183_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17045_ _09569_ _09585_ vssd1 vssd1 vccd1 vccd1 _09586_ sky130_fd_sc_hd__and2_1
XFILLER_171_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14257_ _06914_ _06934_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__nand2_1
X_11469_ rbzero.tex_r1\[2\] _03961_ _03929_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__a21o_1
XFILLER_87_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13208_ _05895_ _05896_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14188_ _06843_ _06876_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__nor2_1
XFILLER_152_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13139_ _05712_ _05718_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__xor2_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18996_ _02658_ vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__clkbuf_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17947_ _01705_ _01707_ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__or2_1
XFILLER_113_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17878_ _01659_ _01660_ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16829_ _09112_ _09116_ _09370_ vssd1 vssd1 vccd1 vccd1 _09371_ sky130_fd_sc_hd__o21ai_1
X_19617_ rbzero.debug_overlay.playerX\[1\] _02982_ rbzero.debug_overlay.playerX\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__o21a_1
XFILLER_96_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19548_ rbzero.pov.spi_buffer\[69\] rbzero.pov.spi_buffer\[70\] _02865_ vssd1 vssd1
+ vccd1 vccd1 _02943_ sky130_fd_sc_hd__mux2_1
XFILLER_59_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19479_ rbzero.pov.spi_buffer\[36\] rbzero.pov.spi_buffer\[37\] _02899_ vssd1 vssd1
+ vccd1 vccd1 _02907_ sky130_fd_sc_hd__mux2_1
XFILLER_62_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21372_ _00395_ _01388_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20323_ gpout0.clk_div\[0\] _03003_ vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__nor2_1
XFILLER_200_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20254_ _03254_ vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__clkinv_2
XFILLER_89_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20185_ _03205_ _03206_ _03207_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__and3_1
XFILLER_77_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10840_ rbzero.tex_g0\[12\] rbzero.tex_g0\[11\] _03638_ vssd1 vssd1 vccd1 vccd1 _03645_
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10771_ rbzero.tex_g0\[45\] rbzero.tex_g0\[44\] _03605_ vssd1 vssd1 vccd1 vccd1 _03609_
+ sky130_fd_sc_hd__mux2_1
XFILLER_198_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12510_ _03789_ _05196_ _05197_ _05198_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_197_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13490_ _05876_ _05874_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__or2b_1
XFILLER_160_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12441_ rbzero.map_rom.a6 _05114_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__or2_1
XFILLER_205_1262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15160_ _07403_ _07751_ _07424_ _07402_ vssd1 vssd1 vccd1 vccd1 _07774_ sky130_fd_sc_hd__o31a_1
XFILLER_172_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12372_ _05056_ _05058_ _05060_ _05063_ _05064_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__a2111o_1
XFILLER_138_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14111_ _05740_ _06423_ _06321_ _06028_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__a2bb2o_1
X_11323_ rbzero.row_render.size\[1\] rbzero.row_render.size\[0\] vssd1 vssd1 vccd1
+ vccd1 _04042_ sky130_fd_sc_hd__nor2_1
XFILLER_197_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15091_ _07341_ _05215_ vssd1 vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__nand2_1
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14042_ _06709_ _06729_ _06730_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__a21oi_1
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11254_ _03968_ _03969_ _03970_ _03971_ _03972_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__o221a_1
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10205_ _03309_ vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_238_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18850_ rbzero.debug_overlay.vplaneY\[-1\] _02541_ vssd1 vssd1 vccd1 vccd1 _02567_
+ sky130_fd_sc_hd__nor2_1
XTAP_6430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11185_ _03903_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__buf_4
XTAP_6441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17801_ _09182_ _09976_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__nor2_1
XTAP_6452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18781_ _02479_ _02491_ _02495_ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__a21oi_1
XTAP_6485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15993_ _07469_ _07805_ vssd1 vssd1 vccd1 vccd1 _08606_ sky130_fd_sc_hd__or2_1
XTAP_5740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17732_ _01447_ _10162_ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__or2b_1
XTAP_5762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14944_ _07498_ _07557_ vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__and2_1
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17663_ _10162_ _01447_ vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__xnor2_1
XFILLER_224_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14875_ _07475_ _07426_ vssd1 vssd1 vccd1 vccd1 _07489_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19402_ rbzero.pov.mosi rbzero.pov.spi_buffer\[0\] _02866_ vssd1 vssd1 vccd1 vccd1
+ _02867_ sky130_fd_sc_hd__mux2_1
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16614_ _09159_ _09222_ vssd1 vssd1 vccd1 vccd1 _09223_ sky130_fd_sc_hd__xnor2_1
XFILLER_211_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13826_ _05668_ _06305_ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__and2_1
X_17594_ _09973_ _09998_ _09997_ vssd1 vssd1 vccd1 vccd1 _10131_ sky130_fd_sc_hd__a21boi_1
XFILLER_235_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19333_ _02856_ vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__clkinv_2
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16545_ _09152_ _09153_ vssd1 vssd1 vccd1 vccd1 _09154_ sky130_fd_sc_hd__nor2_1
XFILLER_1_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13757_ _06432_ _06445_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__nor2_1
XFILLER_188_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10969_ _03712_ vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12708_ _05361_ _05363_ _05376_ _05396_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__or4_2
X_19264_ _02816_ vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__clkbuf_1
XFILLER_231_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16476_ _08881_ _08948_ _09085_ vssd1 vssd1 vccd1 vccd1 _09086_ sky130_fd_sc_hd__a21bo_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13688_ _06327_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__inv_2
X_18215_ _01990_ _01994_ rbzero.wall_tracer.trackDistX\[11\] _09276_ vssd1 vssd1 vccd1
+ vccd1 _00564_ sky130_fd_sc_hd__o2bb2a_1
X_15427_ _07443_ _07709_ _08038_ vssd1 vssd1 vccd1 vccd1 _08041_ sky130_fd_sc_hd__or3_1
XFILLER_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12639_ _05325_ _05327_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__or2_1
XFILLER_54_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19195_ rbzero.spi_registers.new_vshift\[1\] _02775_ vssd1 vssd1 vccd1 vccd1 _02777_
+ sky130_fd_sc_hd__or2_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18146_ _08595_ _09051_ vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__nor2_1
XFILLER_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15358_ _07670_ _07971_ vssd1 vssd1 vccd1 vccd1 _07972_ sky130_fd_sc_hd__or2_1
XFILLER_129_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14309_ _06573_ _06629_ vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__or2_1
XFILLER_176_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18077_ _09833_ _09373_ _01761_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__or3_1
XFILLER_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15289_ _07875_ _07902_ vssd1 vssd1 vccd1 vccd1 _07903_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17028_ _09448_ _09458_ _09457_ vssd1 vssd1 vccd1 vccd1 _09569_ sky130_fd_sc_hd__a21bo_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18979_ _02649_ vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__clkbuf_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20941_ net104 _00957_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20872_ net59 _00888_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21355_ _00378_ _01371_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20306_ _02855_ vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__clkinv_2
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21286_ _00335_ _01302_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20237_ _03246_ _03249_ _03250_ _09244_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__a31o_1
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20168_ rbzero.traced_texa\[0\] rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1 _03194_
+ sky130_fd_sc_hd__nand2_1
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12990_ _05626_ _05630_ _05591_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__a21oi_1
X_20099_ _02708_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__clkbuf_4
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11941_ _04611_ _04618_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__nor2_1
XFILLER_233_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14660_ _03800_ _07302_ _07303_ _07257_ vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__o211a_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _03984_ _04577_ _04585_ _04026_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__a31o_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _06291_ _06299_ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__xnor2_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10823_ rbzero.tex_g0\[20\] rbzero.tex_g0\[19\] _03627_ vssd1 vssd1 vccd1 vccd1 _03636_
+ sky130_fd_sc_hd__mux2_1
XFILLER_207_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14591_ _05018_ _07254_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__nor2_1
XFILLER_26_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16330_ _08914_ _08940_ vssd1 vssd1 vccd1 vccd1 _08941_ sky130_fd_sc_hd__xor2_1
XFILLER_38_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13542_ _06230_ _05848_ vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__nand2_1
XFILLER_213_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10754_ _03599_ vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16261_ _08737_ _08730_ vssd1 vssd1 vccd1 vccd1 _08872_ sky130_fd_sc_hd__and2b_1
XFILLER_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13473_ _05934_ _05980_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__nor2_1
XFILLER_16_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10685_ rbzero.tex_g1\[21\] rbzero.tex_g1\[22\] _03563_ vssd1 vssd1 vccd1 vccd1 _03564_
+ sky130_fd_sc_hd__mux2_1
X_18000_ _08732_ _08645_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__nor2_1
XFILLER_200_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15212_ _07470_ vssd1 vssd1 vccd1 vccd1 _07826_ sky130_fd_sc_hd__buf_4
XFILLER_142_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12424_ _05115_ _05116_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__nor2_1
XFILLER_127_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16192_ _08639_ _08649_ _08803_ vssd1 vssd1 vccd1 vccd1 _08804_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15143_ _07724_ _07738_ vssd1 vssd1 vccd1 vccd1 _07757_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12355_ _05037_ _05043_ _05044_ _05047_ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__and4b_1
XFILLER_86_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11306_ _04007_ _04020_ _04024_ _03899_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__a211o_1
X_15074_ _07217_ _07687_ vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__nor2_1
X_12286_ _04979_ rbzero.wall_tracer.trackDistY\[-5\] _04977_ rbzero.wall_tracer.trackDistY\[-6\]
+ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__a22o_1
XFILLER_138_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19951_ _03118_ vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__clkinv_2
XFILLER_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14025_ _06673_ _06672_ _06664_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__a21o_1
X_18902_ _02609_ vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__clkbuf_1
X_11237_ _03949_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__buf_4
XFILLER_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19882_ _03111_ vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__clkinv_2
XFILLER_214_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11168_ _03879_ _03884_ _03885_ _03886_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__o211a_1
X_18833_ _02538_ _02541_ _02550_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__a21oi_1
XTAP_6260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18764_ _02472_ rbzero.wall_tracer.rayAddendY\[4\] vssd1 vssd1 vccd1 vccd1 _02487_
+ sky130_fd_sc_hd__xnor2_1
XTAP_5570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15976_ _08557_ _08559_ vssd1 vssd1 vccd1 vccd1 _08589_ sky130_fd_sc_hd__or2_1
XFILLER_110_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11099_ _03818_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__buf_4
XFILLER_222_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17715_ _01498_ _01499_ vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__nand2_2
XFILLER_209_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14927_ _07356_ _07540_ vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__nand2_1
XFILLER_110_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18695_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__nand2_1
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17646_ _10096_ _10098_ _10094_ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__a21bo_1
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14858_ _07455_ vssd1 vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__clkbuf_4
XFILLER_184_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13809_ _06458_ _06477_ _06497_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__o21a_1
X_17577_ _07858_ _09603_ _10112_ _10113_ vssd1 vssd1 vccd1 vccd1 _10114_ sky130_fd_sc_hd__or4bb_1
XFILLER_189_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14789_ _07380_ _07401_ _07402_ vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__o21ai_1
XFILLER_205_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19316_ rbzero.pov.spi_counter\[3\] _02846_ _02848_ _02844_ vssd1 vssd1 vccd1 vccd1
+ _00811_ sky130_fd_sc_hd__o211a_1
X_16528_ _09135_ _09136_ vssd1 vssd1 vccd1 vccd1 _09137_ sky130_fd_sc_hd__and2_1
XFILLER_189_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19247_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.new_leak\[2\] _02804_
+ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__mux2_1
X_16459_ _09065_ _09066_ _09068_ vssd1 vssd1 vccd1 vccd1 _09069_ sky130_fd_sc_hd__nand3_1
XFILLER_34_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19178_ rbzero.spi_registers.new_floor\[1\] rbzero.spi_registers.got_new_floor _02724_
+ _02753_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__a31o_1
XFILLER_129_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18129_ _01814_ _01816_ _01909_ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__o21a_1
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21140_ _00189_ _01156_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21071_ _00120_ _01087_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20022_ _03124_ vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__clkinv_2
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20924_ net75 _00940_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20855_ _00073_ _00871_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20786_ net102 _00802_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10470_ rbzero.tex_r0\[60\] rbzero.tex_r0\[59\] _03446_ vssd1 vssd1 vccd1 vccd1 _03451_
+ sky130_fd_sc_hd__mux2_1
XFILLER_202_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21407_ net115 _01423_ vssd1 vssd1 vccd1 vccd1 gpout4.clk_div\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12140_ _04843_ _04845_ _04846_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__and3_1
XFILLER_151_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21338_ _00361_ _01354_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12071_ net24 net23 vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__nor2_1
XFILLER_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21269_ _00318_ _01285_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11022_ _03740_ _03741_ _03747_ _03749_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__a31o_1
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15830_ _08353_ _08354_ _08416_ _08443_ vssd1 vssd1 vccd1 vccd1 _08444_ sky130_fd_sc_hd__o22a_1
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15761_ _08358_ _08359_ _08374_ vssd1 vssd1 vccd1 vccd1 _08375_ sky130_fd_sc_hd__a21o_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ _05433_ _05660_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__or2_1
XFILLER_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17500_ _10014_ _09900_ vssd1 vssd1 vccd1 vccd1 _10037_ sky130_fd_sc_hd__or2b_1
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14712_ _07330_ vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_206_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11924_ _03294_ _03295_ gpout0.vpos\[8\] _04110_ net9 _04625_ vssd1 vssd1 vccd1 vccd1
+ _04635_ sky130_fd_sc_hd__mux4_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ _02226_ _02227_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__nand2_1
X_15692_ _08291_ _08305_ vssd1 vssd1 vccd1 vccd1 _08306_ sky130_fd_sc_hd__xnor2_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17431_ _09968_ _08780_ _09838_ _09837_ vssd1 vssd1 vccd1 vccd1 _09969_ sky130_fd_sc_hd__o31a_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _07291_ _07246_ _07249_ vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__o21ai_1
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _03898_ _04560_ _04568_ _03953_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__o211a_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17362_ _09653_ _09655_ _09787_ _09785_ vssd1 vssd1 vccd1 vccd1 _09900_ sky130_fd_sc_hd__a31o_1
XFILLER_199_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10806_ _03604_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__clkbuf_4
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14574_ _07101_ _07240_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__nand2_1
XFILLER_158_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11786_ _04498_ _04499_ _04500_ _04323_ _03972_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__o221a_1
XFILLER_213_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19101_ _02714_ vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__clkbuf_1
X_16313_ _08917_ _08923_ _07697_ _07698_ vssd1 vssd1 vccd1 vccd1 _08924_ sky130_fd_sc_hd__and4bb_1
XFILLER_198_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13525_ _05872_ _06179_ _06213_ vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__a21oi_2
XFILLER_158_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17293_ _09830_ _09831_ vssd1 vssd1 vccd1 vccd1 _09832_ sky130_fd_sc_hd__nand2_1
XFILLER_144_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10737_ _03590_ vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19032_ _02677_ vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16244_ _04938_ _08663_ vssd1 vssd1 vccd1 vccd1 _08855_ sky130_fd_sc_hd__nor2_2
XFILLER_186_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13456_ _06092_ _06096_ _06121_ _06144_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__and4_1
XFILLER_173_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10668_ rbzero.tex_g1\[29\] rbzero.tex_g1\[30\] _03552_ vssd1 vssd1 vccd1 vccd1 _03555_
+ sky130_fd_sc_hd__mux2_1
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ _05056_ _05099_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__and2_1
X_16175_ _08785_ vssd1 vssd1 vccd1 vccd1 _08787_ sky130_fd_sc_hd__clkbuf_4
X_13387_ _05627_ _05635_ _05657_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__or3_1
X_10599_ _03518_ vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15126_ _07724_ _07738_ _07739_ vssd1 vssd1 vccd1 vccd1 _07740_ sky130_fd_sc_hd__a21oi_1
X_12338_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__nand2_1
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15057_ _03794_ rbzero.wall_tracer.stepDistY\[0\] vssd1 vssd1 vccd1 vccd1 _07671_
+ sky130_fd_sc_hd__nor2_1
XFILLER_138_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19934_ _03116_ vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__clkinv_2
X_12269_ rbzero.wall_tracer.trackDistX\[-8\] vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__inv_2
XFILLER_218_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14008_ _06694_ _06695_ vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19865_ _03109_ vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__clkinv_2
XFILLER_96_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18816_ _02509_ rbzero.debug_overlay.vplaneY\[-1\] vssd1 vssd1 vccd1 vccd1 _02536_
+ sky130_fd_sc_hd__and2_1
XTAP_6090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19796_ _03096_ _03097_ vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__nor2_1
XFILLER_83_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15959_ _08171_ _08457_ vssd1 vssd1 vccd1 vccd1 _08573_ sky130_fd_sc_hd__xnor2_4
X_18747_ _02471_ vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18678_ rbzero.debug_overlay.vplaneY\[-2\] rbzero.wall_tracer.rayAddendY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__or2_1
XFILLER_224_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17629_ _09684_ _08851_ _08979_ _09022_ vssd1 vssd1 vccd1 vccd1 _10165_ sky130_fd_sc_hd__o22a_1
XFILLER_211_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20640_ net56 _00656_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20571_ net125 _00587_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21123_ _00172_ _01139_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21054_ _00103_ _01070_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20005_ _03123_ vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__clkinv_2
XFILLER_189_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ net61 _00923_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[44\] sky130_fd_sc_hd__dfxtp_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ rbzero.tex_g0\[46\] _03925_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__and2_1
X_20838_ _00056_ _00854_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_243_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11571_ rbzero.debug_overlay.playerX\[-5\] _04214_ _04237_ rbzero.debug_overlay.playerX\[-6\]
+ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__a22o_1
XFILLER_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20769_ net103 _00785_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13310_ _05967_ _05998_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__or2_1
XFILLER_168_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10522_ rbzero.tex_r0\[35\] rbzero.tex_r0\[34\] _03468_ vssd1 vssd1 vccd1 vccd1 _03478_
+ sky130_fd_sc_hd__mux2_1
X_14290_ _06371_ _06402_ _06975_ _06978_ vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__o31a_2
XFILLER_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13241_ _05905_ _05929_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__xnor2_1
X_10453_ rbzero.tex_r1\[1\] rbzero.tex_r1\[2\] _03433_ vssd1 vssd1 vccd1 vccd1 _03440_
+ sky130_fd_sc_hd__mux2_1
XFILLER_164_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13172_ _05401_ _05703_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__nand2_4
X_10384_ rbzero.tex_r1\[34\] rbzero.tex_r1\[35\] _03400_ vssd1 vssd1 vccd1 vccd1 _03404_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ net30 net29 vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__nor2_1
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17980_ _09429_ _09373_ _01761_ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__or3_1
XFILLER_215_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16931_ _09471_ _09472_ vssd1 vssd1 vccd1 vccd1 _09473_ sky130_fd_sc_hd__xnor2_1
X_12054_ net49 net40 net39 net41 _04718_ _04717_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__mux4_1
XFILLER_117_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11005_ rbzero.map_rom.b6 vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__buf_2
XFILLER_237_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16862_ _09143_ _09146_ _09145_ vssd1 vssd1 vccd1 vccd1 _09404_ sky130_fd_sc_hd__a21bo_1
X_19650_ _07458_ _02958_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__nor2_1
XFILLER_133_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15813_ _08424_ _08426_ _08418_ vssd1 vssd1 vccd1 vccd1 _08427_ sky130_fd_sc_hd__a21o_1
X_18601_ _02338_ _02339_ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__nor2_1
X_19581_ rbzero.pov.ready_buffer\[60\] _07432_ _02963_ vssd1 vssd1 vccd1 vccd1 _02964_
+ sky130_fd_sc_hd__mux2_1
XFILLER_133_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16793_ rbzero.wall_tracer.trackDistX\[-4\] rbzero.wall_tracer.stepDistX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _09339_ sky130_fd_sc_hd__nor2_1
XFILLER_19_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18532_ rbzero.wall_tracer.rayAddendX\[4\] rbzero.wall_tracer.rayAddendX\[3\] _02275_
+ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__o21ai_1
X_15744_ _08341_ _08339_ _08340_ vssd1 vssd1 vccd1 vccd1 _08358_ sky130_fd_sc_hd__nand3_1
XFILLER_19_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12956_ _05608_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__clkinv_2
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ net10 vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__buf_2
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18463_ _02198_ _02209_ _02210_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__or3_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ _08234_ _08288_ vssd1 vssd1 vccd1 vccd1 _08289_ sky130_fd_sc_hd__and2b_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _05568_ _05570_ _05574_ _05575_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__or4_1
XFILLER_60_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _09835_ _09843_ _09951_ vssd1 vssd1 vccd1 vccd1 _09952_ sky130_fd_sc_hd__a21o_1
XFILLER_206_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ rbzero.wall_tracer.trackDistX\[-1\] rbzero.wall_tracer.trackDistY\[-1\] _07258_
+ vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__mux2_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _03920_ _04547_ _04551_ _03898_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__a211o_1
X_18394_ rbzero.debug_overlay.vplaneX\[-9\] rbzero.wall_tracer.rayAddendX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__nand2_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _09773_ _09774_ _09882_ vssd1 vssd1 vccd1 vccd1 _09884_ sky130_fd_sc_hd__a21o_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14557_ _07029_ _06985_ _05568_ _07031_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__or4b_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11769_ _04482_ _04483_ _03968_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__mux2_1
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13508_ _05862_ _05864_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__and2b_1
X_17276_ _09809_ _09814_ vssd1 vssd1 vccd1 vccd1 _09815_ sky130_fd_sc_hd__nor2_1
XFILLER_147_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14488_ _07102_ _07171_ vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__nand2_2
XFILLER_147_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19015_ _02668_ vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__clkbuf_1
X_16227_ _08832_ _08834_ _08831_ vssd1 vssd1 vccd1 vccd1 _08838_ sky130_fd_sc_hd__o21bai_1
XFILLER_70_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13439_ _06108_ _06109_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__nand2_1
XFILLER_31_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16158_ _08627_ _08637_ _08635_ vssd1 vssd1 vccd1 vccd1 _08770_ sky130_fd_sc_hd__a21boi_1
XFILLER_161_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15109_ _07717_ _07719_ _07722_ vssd1 vssd1 vccd1 vccd1 _07723_ sky130_fd_sc_hd__a21boi_1
XFILLER_177_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16089_ _08700_ _08701_ vssd1 vssd1 vccd1 vccd1 _08702_ sky130_fd_sc_hd__nor2_1
XFILLER_103_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19917_ _03115_ vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__clkinv_2
XFILLER_151_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19848_ _02862_ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__buf_4
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19779_ _04631_ _03808_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__nand2_1
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20623_ net79 _00639_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20554_ net120 _00570_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20485_ net111 _00501_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21106_ _00155_ _01122_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_6837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout120 net122 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_2
XFILLER_134_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout131 net140 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_2
X_21037_ _00086_ _01053_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12810_ _05460_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__buf_2
XFILLER_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13790_ _05767_ _06422_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__or2_1
XFILLER_90_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12741_ _05429_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__clkbuf_4
XFILLER_128_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _08027_ _08029_ vssd1 vssd1 vccd1 vccd1 _08074_ sky130_fd_sc_hd__xnor2_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12672_ _05310_ _05322_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__nand2_2
XFILLER_203_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _07099_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__clkbuf_4
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ rbzero.tex_g0\[55\] rbzero.tex_g0\[54\] _04148_ vssd1 vssd1 vccd1 vccd1 _04340_
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15391_ _07947_ _07948_ vssd1 vssd1 vccd1 vccd1 _08005_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17130_ _09668_ _09669_ vssd1 vssd1 vccd1 vccd1 _09670_ sky130_fd_sc_hd__nand2_1
X_14342_ _06981_ _06980_ _07030_ vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__a21o_1
XFILLER_180_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11554_ rbzero.debug_overlay.facingY\[-6\] _04237_ _04238_ rbzero.debug_overlay.facingY\[-7\]
+ _04271_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__a221o_1
XFILLER_195_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17061_ _08922_ _09470_ vssd1 vssd1 vccd1 vccd1 _09602_ sky130_fd_sc_hd__and2_1
XFILLER_183_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10505_ _03469_ vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__clkbuf_1
X_14273_ _06795_ _06877_ _06879_ _06959_ _06961_ vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__a32o_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11485_ _03823_ _04202_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__nand2_2
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16012_ _08615_ _08623_ vssd1 vssd1 vccd1 vccd1 _08625_ sky130_fd_sc_hd__or2_1
X_13224_ _05672_ _05604_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__nor2_1
XFILLER_143_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10436_ rbzero.tex_r1\[9\] rbzero.tex_r1\[10\] _03422_ vssd1 vssd1 vccd1 vccd1 _03431_
+ sky130_fd_sc_hd__mux2_1
XFILLER_171_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13155_ _05761_ _05779_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__and2_1
XFILLER_87_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10367_ rbzero.tex_r1\[42\] rbzero.tex_r1\[43\] _03389_ vssd1 vssd1 vccd1 vccd1 _03395_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12106_ _04773_ net21 gpout3.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__and3_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17963_ _09968_ _09978_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__nor2_1
XFILLER_215_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13086_ _05769_ _05770_ _05774_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__o21ai_2
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _03358_ vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19702_ _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__buf_2
XFILLER_239_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16914_ _09454_ _09455_ vssd1 vssd1 vccd1 vccd1 _09456_ sky130_fd_sc_hd__xnor2_1
XFILLER_214_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12037_ _04742_ _04744_ _04745_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__and3_1
XFILLER_61_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17894_ _01670_ _01676_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__xnor2_1
XFILLER_239_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19633_ _02999_ _03002_ _03003_ vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__a21oi_1
XFILLER_238_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16845_ _09385_ _09386_ vssd1 vssd1 vccd1 vccd1 _09387_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16776_ _07332_ _08564_ vssd1 vssd1 vccd1 vccd1 _09324_ sky130_fd_sc_hd__and2_1
X_19564_ net53 rbzero.pov.sclk_buffer\[0\] _02708_ vssd1 vssd1 vccd1 vccd1 _02951_
+ sky130_fd_sc_hd__mux2_1
XFILLER_230_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13988_ _06661_ _06675_ _06676_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15727_ _08333_ _08334_ _08338_ vssd1 vssd1 vccd1 vccd1 _08341_ sky130_fd_sc_hd__nand3_1
X_18515_ _02252_ _02253_ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__or2_1
X_12939_ _05467_ _05500_ _05511_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__o21a_1
XFILLER_94_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19495_ _02915_ vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__clkbuf_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15658_ _07379_ vssd1 vssd1 vccd1 vccd1 _08272_ sky130_fd_sc_hd__buf_4
XFILLER_59_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18446_ _02190_ _02192_ _02193_ _02181_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__a22o_1
XFILLER_233_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14609_ _07245_ _07267_ _07268_ _07251_ vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__o211a_1
X_18377_ _02126_ _02132_ _02131_ _09351_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__a31o_1
X_15589_ _08202_ _07842_ vssd1 vssd1 vccd1 vccd1 _08203_ sky130_fd_sc_hd__nor2_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17328_ _09737_ _09738_ vssd1 vssd1 vccd1 vccd1 _09867_ sky130_fd_sc_hd__nor2_1
XFILLER_187_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17259_ _08135_ _08855_ _09797_ vssd1 vssd1 vccd1 vccd1 _09798_ sky130_fd_sc_hd__a21oi_1
XFILLER_147_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20270_ _03255_ vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__clkinv_2
XFILLER_192_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20606_ net90 _00622_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20537_ net136 _00553_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20468_ net119 _00484_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[3\] sky130_fd_sc_hd__dfxtp_1
X_11270_ _03987_ _03988_ _03930_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__mux2_1
XFILLER_197_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10221_ rbzero.tex_b1\[47\] rbzero.tex_b1\[48\] _03311_ vssd1 vssd1 vccd1 vccd1 _03318_
+ sky130_fd_sc_hd__mux2_1
X_20399_ net121 _00430_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_79_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14960_ _07571_ _07572_ _07573_ vssd1 vssd1 vccd1 vccd1 _07574_ sky130_fd_sc_hd__a21o_1
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13911_ _06593_ _06598_ _06599_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__o21a_1
XTAP_5977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14891_ _07502_ _07504_ _07351_ vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__a21o_1
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16630_ _08585_ _09238_ vssd1 vssd1 vccd1 vccd1 _09239_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13842_ _06313_ _06331_ _06526_ _06530_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__o31ai_1
XFILLER_63_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16561_ _07890_ _08636_ vssd1 vssd1 vccd1 vccd1 _09170_ sky130_fd_sc_hd__or2b_1
XFILLER_244_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13773_ _06115_ _06320_ _06461_ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__nand3_1
XFILLER_245_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10985_ rbzero.tex_b0\[7\] rbzero.tex_b0\[6\] _03715_ vssd1 vssd1 vccd1 vccd1 _03721_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18300_ _02066_ _02061_ _02064_ _02065_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__a211oi_2
X_15512_ _08122_ _08124_ _08125_ vssd1 vssd1 vccd1 vccd1 _08126_ sky130_fd_sc_hd__a21boi_1
X_12724_ _05298_ _05412_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__nand2_1
X_19280_ rbzero.spi_registers.spi_cmd\[3\] _02581_ _02578_ rbzero.spi_registers.spi_done
+ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__or4b_1
XFILLER_245_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16492_ _09099_ _09100_ vssd1 vssd1 vccd1 vccd1 _09102_ sky130_fd_sc_hd__nand2_1
XFILLER_200_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18231_ _02004_ _02005_ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__and2_1
X_15443_ _07567_ _07986_ vssd1 vssd1 vccd1 vccd1 _08057_ sky130_fd_sc_hd__nor2_1
XFILLER_54_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12655_ _05343_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__inv_2
XFILLER_54_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18162_ _08781_ _08784_ _08732_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__a21o_1
XFILLER_15_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11606_ _03910_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__buf_4
XFILLER_54_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15374_ _07508_ _07542_ _07550_ _07593_ vssd1 vssd1 vccd1 vccd1 _07988_ sky130_fd_sc_hd__o22ai_1
XFILLER_141_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12586_ _03816_ _05104_ _05105_ _05274_ _03789_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__a311o_1
X_17113_ _09535_ _09544_ _09542_ vssd1 vssd1 vccd1 vccd1 _09653_ sky130_fd_sc_hd__a21o_1
X_14325_ _07012_ _07013_ vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18093_ _07619_ _08634_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__nor2_1
XFILLER_209_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11537_ rbzero.debug_overlay.vplaneX\[-2\] _04245_ _04243_ rbzero.debug_overlay.vplaneX\[0\]
+ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__a221o_1
XFILLER_106_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17044_ _09575_ _09584_ vssd1 vssd1 vccd1 vccd1 _09585_ sky130_fd_sc_hd__xor2_1
XFILLER_183_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14256_ _06799_ _06937_ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__or2_1
XFILLER_176_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11468_ rbzero.tex_r1\[3\] _04142_ _04144_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__and3_1
XFILLER_143_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13207_ _05525_ _05567_ _05748_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__and3_1
X_10419_ _03388_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__clkbuf_4
X_14187_ _06851_ _06874_ _06875_ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__o21ba_1
XFILLER_174_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11399_ _03826_ _04100_ _04117_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__o21bai_4
XFILLER_225_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _05808_ _05812_ _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__a21o_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18995_ rbzero.pov.spi_buffer\[45\] rbzero.pov.ready_buffer\[45\] _02651_ vssd1 vssd1
+ vccd1 vccd1 _02658_ sky130_fd_sc_hd__mux2_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17946_ _01702_ _01704_ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__or2_1
X_13069_ _05756_ _05757_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__or2_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17877_ _07670_ _08723_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__or2_1
XFILLER_113_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19616_ rbzero.debug_overlay.playerX\[1\] _02956_ _02988_ _02989_ vssd1 vssd1 vccd1
+ vccd1 _00970_ sky130_fd_sc_hd__a211o_1
XFILLER_66_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16828_ _09110_ _08989_ _08990_ vssd1 vssd1 vccd1 vccd1 _09370_ sky130_fd_sc_hd__or3_1
XFILLER_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19547_ _02942_ vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__clkbuf_1
X_16759_ rbzero.wall_tracer.trackDistX\[-9\] _09301_ _09302_ _09309_ vssd1 vssd1 vccd1
+ vccd1 _00544_ sky130_fd_sc_hd__o22a_1
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19478_ _02906_ vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18429_ _02180_ vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21371_ _00394_ _01387_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20322_ rbzero.traced_texVinit\[11\] _03260_ _09267_ _09887_ vssd1 vssd1 vccd1 vccd1
+ _01405_ sky130_fd_sc_hd__a22o_1
XFILLER_107_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20253_ _03254_ vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__clkinv_2
XFILLER_66_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20184_ _03205_ _03206_ _03207_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__a21o_1
XFILLER_130_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10770_ _03608_ vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12440_ rbzero.map_rom.a6 _05114_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__nand2_1
XFILLER_51_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12371_ rbzero.debug_overlay.facingY\[0\] rbzero.wall_tracer.rayAddendY\[8\] vssd1
+ vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__nor2_1
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14110_ _06137_ _06423_ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__nor2_1
XFILLER_166_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11322_ rbzero.row_render.size\[2\] vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__inv_2
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15090_ _07444_ _07703_ _07337_ vssd1 vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__a21o_1
XFILLER_180_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14041_ _06710_ _06728_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__and2b_1
XFILLER_84_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11253_ _03945_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__buf_4
XTAP_7121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10204_ rbzero.tex_b1\[55\] rbzero.tex_b1\[56\] _03300_ vssd1 vssd1 vccd1 vccd1 _03309_
+ sky130_fd_sc_hd__mux2_1
XTAP_6420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11184_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__buf_2
XTAP_6431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17800_ _01472_ _01474_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__nand2_1
XTAP_6453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15992_ _08602_ _08604_ vssd1 vssd1 vccd1 vccd1 _08605_ sky130_fd_sc_hd__nand2_1
XFILLER_0_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18780_ _02500_ _02501_ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__nor2_1
XTAP_6475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17731_ _10041_ _10160_ _10158_ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__a21o_1
XTAP_5763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14943_ rbzero.debug_overlay.playerY\[-2\] _07497_ rbzero.debug_overlay.playerY\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _07557_ sky130_fd_sc_hd__o21ai_1
XFILLER_248_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17662_ _01445_ _01446_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__nand2_1
X_14874_ _07477_ _07486_ _07487_ vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__a21bo_1
XFILLER_1_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19401_ _02865_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__clkbuf_4
X_16613_ _09220_ _09221_ vssd1 vssd1 vccd1 vccd1 _09222_ sky130_fd_sc_hd__xor2_1
X_13825_ _05668_ _06311_ _06513_ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__a21o_1
X_17593_ _10128_ _10129_ vssd1 vssd1 vccd1 vccd1 _10130_ sky130_fd_sc_hd__or2_1
XFILLER_169_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16544_ _09149_ _09151_ vssd1 vssd1 vccd1 vccd1 _09153_ sky130_fd_sc_hd__and2_1
X_19332_ _02856_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__clkinv_2
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13756_ _06434_ _06443_ _06444_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__a21boi_1
XFILLER_204_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10968_ rbzero.tex_b0\[15\] rbzero.tex_b0\[14\] _03704_ vssd1 vssd1 vccd1 vccd1 _03712_
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12707_ _05394_ _05378_ _05381_ _05395_ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__or4_1
X_16475_ _08945_ _08947_ vssd1 vssd1 vccd1 vccd1 _09085_ sky130_fd_sc_hd__nand2_1
XFILLER_189_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19263_ rbzero.spi_registers.new_other\[2\] rbzero.spi_registers.spi_buffer\[2\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__mux2_1
XFILLER_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13687_ _06328_ _06375_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__nand2_1
X_10899_ rbzero.tex_b0\[48\] rbzero.tex_b0\[47\] _03671_ vssd1 vssd1 vccd1 vccd1 _03676_
+ sky130_fd_sc_hd__mux2_1
X_18214_ _07332_ _01993_ _09275_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__o21a_1
XFILLER_188_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15426_ _08038_ _08039_ vssd1 vssd1 vccd1 vccd1 _08040_ sky130_fd_sc_hd__xnor2_1
X_12638_ _05276_ _05326_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__xnor2_2
X_19194_ rbzero.spi_registers.vshift\[0\] _02774_ _02776_ _02738_ vssd1 vssd1 vccd1
+ vccd1 _00761_ sky130_fd_sc_hd__o211a_1
XFILLER_141_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18145_ _01861_ _01870_ _01868_ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__a21o_1
X_15357_ _07970_ vssd1 vssd1 vccd1 vccd1 _07971_ sky130_fd_sc_hd__clkbuf_4
XFILLER_200_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12569_ _05149_ _05257_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__and2_1
XFILLER_184_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14308_ _05431_ _06996_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__and2_1
XFILLER_184_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18076_ _09833_ _08852_ _09373_ _07760_ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__o22a_1
XFILLER_184_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15288_ _07900_ _07901_ vssd1 vssd1 vccd1 vccd1 _07902_ sky130_fd_sc_hd__nand2_1
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17027_ _09433_ _09441_ _09567_ vssd1 vssd1 vccd1 vccd1 _09568_ sky130_fd_sc_hd__a21o_1
X_14239_ _06911_ _06926_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__nand2_1
XFILLER_217_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18978_ rbzero.pov.spi_buffer\[37\] rbzero.pov.ready_buffer\[37\] _02640_ vssd1 vssd1
+ vccd1 vccd1 _02649_ sky130_fd_sc_hd__mux2_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _01708_ _01710_ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__nand2_1
XFILLER_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20940_ net85 _00956_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ss_buffer\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20871_ net54 _00887_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21354_ _00377_ _01370_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20305_ _02855_ vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__clkinv_2
XFILLER_194_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21285_ _00334_ _01301_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20236_ _03246_ _03249_ _03250_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__a21oi_1
XFILLER_235_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20167_ rbzero.traced_texa\[0\] rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1 _03193_
+ sky130_fd_sc_hd__or2_1
XFILLER_104_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20098_ rbzero.traced_texa\[-12\] rbzero.texV\[-12\] vssd1 vssd1 vccd1 vccd1 _03136_
+ sky130_fd_sc_hd__or2_1
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ net13 net14 vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__and2b_1
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11871_ _03920_ _04580_ _04584_ _03898_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__a211o_1
XFILLER_79_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13610_ _06292_ _06298_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10822_ _03635_ vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _05025_ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__inv_2
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13541_ _05610_ vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__inv_2
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10753_ rbzero.tex_g0\[53\] rbzero.tex_g0\[52\] _03593_ vssd1 vssd1 vccd1 vccd1 _03599_
+ sky130_fd_sc_hd__mux2_1
XFILLER_207_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16260_ _08863_ _08870_ vssd1 vssd1 vccd1 vccd1 _08871_ sky130_fd_sc_hd__xnor2_1
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ _05979_ _06025_ _06158_ _06160_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__a22o_1
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10684_ _03388_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__clkbuf_4
XFILLER_51_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15211_ _07470_ _07471_ _07817_ _07824_ vssd1 vssd1 vccd1 vccd1 _07825_ sky130_fd_sc_hd__or4_1
XFILLER_16_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12423_ rbzero.map_rom.c6 _05114_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__nor2_1
XFILLER_127_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16191_ _08647_ _08648_ vssd1 vssd1 vccd1 vccd1 _08803_ sky130_fd_sc_hd__nor2_1
XFILLER_200_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15142_ _07741_ _07755_ vssd1 vssd1 vccd1 vccd1 _07756_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12354_ _05045_ _05046_ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__and2_1
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11305_ _04021_ _04022_ _04023_ _03932_ _03946_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__o221a_1
X_15073_ _07202_ _07444_ _07211_ _07208_ _07206_ vssd1 vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__a2111o_1
XFILLER_5_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19950_ _03118_ vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__clkinv_2
X_12285_ rbzero.wall_tracer.trackDistX\[-5\] vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__inv_2
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14024_ _06673_ _06664_ _06672_ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__nand3_1
X_18901_ rbzero.pov.spi_buffer\[0\] rbzero.pov.ready_buffer\[0\] _02608_ vssd1 vssd1
+ vccd1 vccd1 _02609_ sky130_fd_sc_hd__mux2_1
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11236_ _03900_ _03922_ _03951_ _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__o211a_1
X_19881_ _02862_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__buf_4
XFILLER_218_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18832_ _02538_ _02541_ _02550_ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__and3_1
XTAP_6250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11167_ _03882_ _03883_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__nand2_1
XTAP_6261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18763_ _02287_ _02477_ _02478_ _02486_ vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__a31o_1
XTAP_5560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15975_ _08459_ _08563_ _08561_ vssd1 vssd1 vccd1 vccd1 _08588_ sky130_fd_sc_hd__a21boi_2
XFILLER_114_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11098_ _03801_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__clkbuf_4
XTAP_5571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17714_ _10150_ _10151_ _01497_ vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__nand3_1
XFILLER_222_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14926_ _07537_ _07539_ _07374_ vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__mux2_1
XFILLER_114_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18694_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__or2_1
XFILLER_97_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17645_ _10073_ _10074_ _10076_ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__a21bo_1
XFILLER_75_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14857_ _07443_ vssd1 vssd1 vccd1 vccd1 _07471_ sky130_fd_sc_hd__buf_2
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ _06495_ _06496_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__nand2_1
XFILLER_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17576_ _08272_ _09449_ _09978_ _09976_ vssd1 vssd1 vccd1 vccd1 _10113_ sky130_fd_sc_hd__or4_1
X_14788_ _07355_ _07378_ _07387_ _07399_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__or4_1
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19315_ rbzero.pov.spi_counter\[3\] _02846_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__nand2_1
XFILLER_232_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16527_ _09133_ _09134_ vssd1 vssd1 vccd1 vccd1 _09136_ sky130_fd_sc_hd__nand2_1
X_13739_ _06425_ _06426_ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__nand2_1
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19246_ _02806_ vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__clkbuf_1
X_16458_ _08927_ _08936_ _09067_ vssd1 vssd1 vccd1 vccd1 _09068_ sky130_fd_sc_hd__a21o_1
XFILLER_188_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15409_ _08005_ _08022_ vssd1 vssd1 vccd1 vccd1 _08023_ sky130_fd_sc_hd__xor2_1
X_16389_ _08274_ _08592_ _07620_ _08671_ vssd1 vssd1 vccd1 vccd1 _08999_ sky130_fd_sc_hd__or4_1
X_19177_ _02765_ vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18128_ _01812_ _01813_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__or2_1
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18059_ _01838_ _01839_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__nor2_1
XFILLER_144_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21070_ _00119_ _01086_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20021_ _03124_ vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__clkinv_2
XFILLER_154_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20923_ net74 _00939_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20854_ _00072_ _00870_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20785_ net101 _00801_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21406_ net115 _01422_ vssd1 vssd1 vccd1 vccd1 gpout4.clk_div\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21337_ _00360_ _01353_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12070_ net24 _04770_ _04774_ _04777_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__o211a_1
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21268_ _00317_ _01284_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11021_ _03738_ _03748_ rbzero.map_rom.d6 rbzero.map_rom.c6 vssd1 vssd1 vccd1 vccd1
+ _03749_ sky130_fd_sc_hd__a211oi_1
X_20219_ rbzero.traced_texa\[7\] rbzero.texV\[7\] _03232_ vssd1 vssd1 vccd1 vccd1
+ _03237_ sky130_fd_sc_hd__a21o_1
XFILLER_172_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21199_ _00248_ _01215_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ _08364_ _08372_ _08373_ vssd1 vssd1 vccd1 vccd1 _08374_ sky130_fd_sc_hd__a21o_1
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12972_ _05633_ _05639_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__xnor2_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14711_ rbzero.wall_tracer.stepDistX\[10\] _07241_ _04931_ vssd1 vssd1 vccd1 vccd1
+ _07330_ sky130_fd_sc_hd__mux2_1
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11923_ _04630_ _04633_ _04618_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__o21ba_1
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15691_ _08300_ _08303_ _08304_ vssd1 vssd1 vccd1 vccd1 _08305_ sky130_fd_sc_hd__a21o_1
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ _08760_ vssd1 vssd1 vccd1 vccd1 _09968_ sky130_fd_sc_hd__buf_2
X_14642_ rbzero.wall_tracer.trackDistX\[4\] vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__inv_2
XFILLER_166_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11854_ _03945_ _04563_ _04567_ _03949_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__a211o_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10805_ _03626_ vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__clkbuf_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17361_ _09895_ _09896_ _09897_ vssd1 vssd1 vccd1 vccd1 _09899_ sky130_fd_sc_hd__o21a_1
X_14573_ _05416_ _05408_ _07239_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__or3_1
XFILLER_198_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11785_ rbzero.tex_b0\[1\] rbzero.tex_b0\[0\] _04001_ vssd1 vssd1 vccd1 vccd1 _04500_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19100_ rbzero.spi_registers.sclk_buffer\[1\] rbzero.spi_registers.sclk_buffer\[0\]
+ _09243_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__mux2_1
X_16312_ _08922_ vssd1 vssd1 vccd1 vccd1 _08923_ sky130_fd_sc_hd__clkbuf_4
X_13524_ _06210_ _06212_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__xor2_1
X_17292_ _07520_ _07651_ _08636_ _09163_ vssd1 vssd1 vccd1 vccd1 _09831_ sky130_fd_sc_hd__a22o_1
XFILLER_207_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10736_ rbzero.tex_g0\[61\] rbzero.tex_g0\[60\] _03512_ vssd1 vssd1 vccd1 vccd1 _03590_
+ sky130_fd_sc_hd__mux2_1
XFILLER_198_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16243_ _07792_ _07788_ _08717_ rbzero.wall_tracer.visualWallDist\[7\] vssd1 vssd1
+ vccd1 vccd1 _08854_ sky130_fd_sc_hd__or4b_1
XFILLER_186_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19031_ rbzero.pov.spi_buffer\[62\] rbzero.pov.ready_buffer\[62\] _02673_ vssd1 vssd1
+ vccd1 vccd1 _02677_ sky130_fd_sc_hd__mux2_1
XFILLER_173_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13455_ _06116_ _06117_ _06120_ _06142_ _06143_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__o221ai_1
XFILLER_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ _03554_ vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__clkbuf_1
X_12406_ _05055_ _05048_ _05052_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__or3_1
X_16174_ _07826_ _07471_ _08780_ _08785_ vssd1 vssd1 vccd1 vccd1 _08786_ sky130_fd_sc_hd__or4_1
XFILLER_51_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13386_ _06043_ _06046_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10598_ rbzero.tex_g1\[62\] rbzero.tex_g1\[63\] _03433_ vssd1 vssd1 vccd1 vccd1 _03518_
+ sky130_fd_sc_hd__mux2_1
XFILLER_115_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15125_ _07716_ _07723_ vssd1 vssd1 vccd1 vccd1 _07739_ sky130_fd_sc_hd__nor2_1
XFILLER_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12337_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] vssd1
+ vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__xnor2_2
XFILLER_126_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15056_ _07337_ _07667_ _07669_ vssd1 vssd1 vccd1 vccd1 _07670_ sky130_fd_sc_hd__o21ai_4
X_19933_ _03116_ vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__clkinv_2
X_12268_ rbzero.wall_tracer.trackDistX\[-7\] vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__inv_2
XFILLER_99_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14007_ _06694_ _06695_ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__nand2_1
XFILLER_218_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11219_ _03859_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__clkbuf_4
XFILLER_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19864_ _03109_ vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__clkinv_2
XFILLER_190_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12199_ _04873_ _04874_ _04116_ _04904_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__a31o_1
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18815_ _02509_ rbzero.debug_overlay.vplaneY\[-1\] vssd1 vssd1 vccd1 vccd1 _02535_
+ sky130_fd_sc_hd__nor2_1
XTAP_6080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19795_ _04104_ _03094_ _02742_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__o21ai_1
XFILLER_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18746_ rbzero.wall_tracer.rayAddendY\[2\] _02470_ _03811_ vssd1 vssd1 vccd1 vccd1
+ _02471_ sky130_fd_sc_hd__mux2_1
XTAP_5390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15958_ rbzero.debug_overlay.playerY\[-7\] rbzero.debug_overlay.playerX\[-7\] _07343_
+ vssd1 vssd1 vccd1 vccd1 _08572_ sky130_fd_sc_hd__mux2_1
XFILLER_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14909_ _07518_ _07522_ vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__nand2_1
XFILLER_37_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18677_ _02406_ vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__clkbuf_1
X_15889_ _07888_ _07897_ _07896_ vssd1 vssd1 vccd1 vccd1 _08503_ sky130_fd_sc_hd__a21o_1
XFILLER_184_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17628_ _10108_ _10092_ vssd1 vssd1 vccd1 vccd1 _10164_ sky130_fd_sc_hd__or2b_1
XFILLER_64_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17559_ _08595_ _10095_ _08917_ _08594_ vssd1 vssd1 vccd1 vccd1 _10096_ sky130_fd_sc_hd__o22ai_1
XFILLER_189_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20570_ net125 _00586_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19229_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.new_floor\[1\]
+ _02795_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__mux2_1
XFILLER_176_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21122_ _00171_ _01138_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21053_ _00102_ _01069_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20004_ _03123_ vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__clkinv_2
XFILLER_247_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20906_ net61 _00922_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[43\] sky130_fd_sc_hd__dfxtp_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20837_ _00055_ _00853_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11570_ rbzero.debug_overlay.playerY\[-9\] _04240_ _04277_ _04287_ vssd1 vssd1 vccd1
+ vccd1 _04288_ sky130_fd_sc_hd__a211o_1
X_20768_ net100 _00784_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10521_ _03477_ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20699_ net101 _00715_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13240_ _05925_ _05927_ _05928_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__a21oi_1
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10452_ _03439_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13171_ _05766_ _05701_ _05773_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__and3_1
XFILLER_108_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10383_ _03403_ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12122_ net30 _04822_ _04826_ _04828_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__o211a_1
XFILLER_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16930_ _08335_ _09051_ vssd1 vssd1 vccd1 vccd1 _09472_ sky130_fd_sc_hd__nor2_1
XFILLER_172_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12053_ net43 _04748_ _04749_ _04116_ _04761_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__a221o_1
XFILLER_117_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11004_ rbzero.map_rom.i_row\[4\] vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__inv_2
XFILLER_238_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16861_ _09401_ _09402_ vssd1 vssd1 vccd1 vccd1 _09403_ sky130_fd_sc_hd__nand2_1
XFILLER_42_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18600_ _02327_ _02330_ _02337_ _09269_ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__a31o_1
XFILLER_24_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15812_ _07878_ _08398_ _08425_ vssd1 vssd1 vccd1 vccd1 _08426_ sky130_fd_sc_hd__or3_1
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19580_ _02962_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__clkbuf_4
X_16792_ _09279_ _08828_ vssd1 vssd1 vccd1 vccd1 _09338_ sky130_fd_sc_hd__nor2_1
XFILLER_93_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18531_ _02274_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__clkbuf_4
X_15743_ _08343_ _08345_ vssd1 vssd1 vccd1 vccd1 _08357_ sky130_fd_sc_hd__xnor2_1
X_12955_ _05633_ _05639_ _05643_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__a21o_1
XFILLER_111_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11906_ _04611_ o_rgb[23] _04615_ _04616_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__a211o_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18462_ _02209_ _02210_ _02198_ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__o21ai_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _07379_ _08060_ vssd1 vssd1 vccd1 vccd1 _08288_ sky130_fd_sc_hd__nor2_1
X_12886_ _05406_ _05548_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__nor2_1
XFILLER_34_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _09840_ _09842_ vssd1 vssd1 vccd1 vccd1 _09951_ sky130_fd_sc_hd__nor2_1
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14625_ rbzero.wall_tracer.visualWallDist\[-2\] _07253_ _07278_ _07279_ _07266_ vssd1
+ vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__o221a_1
XFILLER_57_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11837_ _03908_ _04548_ _04549_ _04550_ _03944_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__o221a_1
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18393_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.wall_tracer.rayAddendX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__nand2_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17344_ _09773_ _09774_ _09882_ vssd1 vssd1 vccd1 vccd1 _09883_ sky130_fd_sc_hd__and3_1
X_14556_ _07226_ vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11768_ rbzero.tex_b0\[25\] rbzero.tex_b0\[24\] _04001_ vssd1 vssd1 vccd1 vccd1 _04483_
+ sky130_fd_sc_hd__mux2_1
XFILLER_202_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13507_ _05692_ _05722_ _05772_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__and3_1
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10719_ _03581_ vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__clkbuf_1
X_17275_ _09812_ _09813_ vssd1 vssd1 vccd1 vccd1 _09814_ sky130_fd_sc_hd__xor2_1
X_14487_ _07159_ _07072_ _07168_ _07170_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__o22a_2
XFILLER_158_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11699_ rbzero.tex_g1\[59\] _03964_ _03965_ _03997_ vssd1 vssd1 vccd1 vccd1 _04415_
+ sky130_fd_sc_hd__a31o_1
XFILLER_228_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19014_ rbzero.pov.spi_buffer\[54\] rbzero.pov.ready_buffer\[54\] _02662_ vssd1 vssd1
+ vccd1 vccd1 _02668_ sky130_fd_sc_hd__mux2_1
XFILLER_70_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13438_ _06007_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__inv_2
X_16226_ rbzero.wall_tracer.texu\[2\] _07338_ _07266_ _08837_ vssd1 vssd1 vccd1 vccd1
+ _00483_ sky130_fd_sc_hd__o211a_1
XFILLER_127_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16157_ _08463_ _08617_ _08768_ _08621_ vssd1 vssd1 vccd1 vccd1 _08769_ sky130_fd_sc_hd__a22o_1
X_13369_ _06056_ _06038_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__and2b_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15108_ _07720_ _07721_ vssd1 vssd1 vccd1 vccd1 _07722_ sky130_fd_sc_hd__nand2_1
XFILLER_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16088_ _07389_ _07394_ _07343_ vssd1 vssd1 vccd1 vccd1 _08701_ sky130_fd_sc_hd__mux2_1
XFILLER_9_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15039_ _04928_ _07651_ _07652_ vssd1 vssd1 vccd1 vccd1 _07653_ sky130_fd_sc_hd__and3_1
XFILLER_69_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19916_ _03115_ vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__clkinv_2
XFILLER_111_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19847_ _03107_ vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__clkinv_2
XFILLER_29_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19778_ _03813_ _03084_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__nor2_1
XFILLER_231_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18729_ _02287_ _02446_ _02447_ _02454_ vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__a31o_1
XFILLER_209_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20622_ net80 _00638_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20553_ net120 _00569_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20484_ net111 _00500_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21105_ _00154_ _01121_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout110 net115 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_2
XTAP_6849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout121 net122 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__buf_2
Xfanout132 net133 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21036_ _00085_ _01052_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12740_ _05428_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__clkbuf_4
XFILLER_16_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12671_ _05348_ _05356_ _05359_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__nor3_2
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14410_ _07076_ _07098_ _05538_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__a21o_2
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11622_ _04337_ _04338_ _03909_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__mux2_1
XFILLER_187_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15390_ _07951_ _07952_ vssd1 vssd1 vccd1 vccd1 _08004_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14341_ _06981_ _06368_ _06979_ vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__nor3_2
XFILLER_168_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11553_ rbzero.debug_overlay.facingY\[-5\] _04214_ _04244_ rbzero.debug_overlay.facingY\[-1\]
+ _04270_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__a221o_1
XFILLER_11_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17060_ _09590_ _09600_ vssd1 vssd1 vccd1 vccd1 _09601_ sky130_fd_sc_hd__xor2_1
XFILLER_183_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10504_ rbzero.tex_r0\[44\] rbzero.tex_r0\[43\] _03468_ vssd1 vssd1 vccd1 vccd1 _03469_
+ sky130_fd_sc_hd__mux2_1
X_14272_ _06795_ _06960_ vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__xnor2_2
XFILLER_184_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11484_ _03783_ gpout0.hpos\[5\] _03806_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__nand3_1
XFILLER_184_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16011_ _08615_ _08623_ vssd1 vssd1 vccd1 vccd1 _08624_ sky130_fd_sc_hd__nand2_1
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13223_ _05611_ _05660_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__nor2_1
XFILLER_171_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10435_ _03430_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13154_ _05758_ _05760_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__and2b_1
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10366_ _03394_ vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12105_ _04803_ _04810_ _04812_ _04809_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__a22o_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _01637_ _01743_ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__nand2_1
X_13085_ _05771_ _05773_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10297_ rbzero.tex_b1\[11\] rbzero.tex_b1\[12\] _03355_ vssd1 vssd1 vccd1 vccd1 _03358_
+ sky130_fd_sc_hd__mux2_1
XFILLER_97_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19701_ rbzero.pov.ready _02721_ _02833_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__nand3_2
X_16913_ _07858_ _08780_ vssd1 vssd1 vccd1 vccd1 _09455_ sky130_fd_sc_hd__nor2_1
X_12036_ net6 net7 _04743_ net8 vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__o22a_1
XFILLER_111_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17893_ _01674_ _01675_ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__nand2_1
XFILLER_78_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19632_ _02753_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__buf_4
X_16844_ _07515_ _08978_ vssd1 vssd1 vccd1 vccd1 _09386_ sky130_fd_sc_hd__nor2_1
XFILLER_66_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19563_ _02950_ vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__clkbuf_1
X_16775_ rbzero.wall_tracer.trackDistX\[-7\] _09301_ _09317_ _09323_ vssd1 vssd1 vccd1
+ vccd1 _00546_ sky130_fd_sc_hd__o22a_1
XFILLER_4_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13987_ _06662_ _06674_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__and2b_1
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18514_ _02248_ _02250_ _02257_ _09256_ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__a31o_1
X_15726_ _08325_ _08327_ vssd1 vssd1 vccd1 vccd1 _08340_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12938_ _05471_ _05474_ _05488_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__a21oi_4
X_19494_ rbzero.pov.spi_buffer\[43\] rbzero.pov.spi_buffer\[44\] _02910_ vssd1 vssd1
+ vccd1 vccd1 _02915_ sky130_fd_sc_hd__mux2_1
XFILLER_59_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18445_ _02194_ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__inv_2
X_15657_ _08244_ _08270_ vssd1 vssd1 vccd1 vccd1 _08271_ sky130_fd_sc_hd__xnor2_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _05499_ _05519_ _05557_ _05481_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__a211o_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14608_ rbzero.wall_tracer.visualWallDist\[-7\] _07249_ vssd1 vssd1 vccd1 vccd1 _07268_
+ sky130_fd_sc_hd__or2_1
XFILLER_61_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18376_ _02126_ _02131_ _02132_ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__a21oi_1
X_15588_ _07384_ _07385_ vssd1 vssd1 vccd1 vccd1 _08202_ sky130_fd_sc_hd__and2_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17327_ _09856_ _09865_ vssd1 vssd1 vccd1 vccd1 _09866_ sky130_fd_sc_hd__xor2_1
XFILLER_147_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14539_ _07212_ vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17258_ _09684_ _08717_ vssd1 vssd1 vccd1 vccd1 _09797_ sky130_fd_sc_hd__nor2_1
XFILLER_128_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16209_ _08661_ _08683_ _08820_ vssd1 vssd1 vccd1 vccd1 _08821_ sky130_fd_sc_hd__a21boi_1
XFILLER_161_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17189_ _09465_ _09466_ _09611_ _09607_ _08779_ vssd1 vssd1 vccd1 vccd1 _09729_ sky130_fd_sc_hd__a32o_1
XFILLER_155_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20605_ net81 _00621_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20536_ net131 _00552_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20467_ net127 _00483_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10220_ _03317_ vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20398_ net125 _00429_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_6602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13910_ _06590_ _06592_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__nand2_1
XFILLER_130_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21019_ net94 _01035_ vssd1 vssd1 vccd1 vccd1 rbzero.vga_sync.vsync sky130_fd_sc_hd__dfxtp_1
XFILLER_48_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14890_ _07334_ _05258_ _07503_ vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__o21ai_1
XTAP_5989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13841_ _06266_ _06389_ _06529_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__or3b_1
XFILLER_169_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16560_ _08241_ _07817_ vssd1 vssd1 vccd1 vccd1 _09169_ sky130_fd_sc_hd__nor2_1
XFILLER_204_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13772_ _06313_ _06330_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__nor2_1
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10984_ _03720_ vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15511_ _07435_ _07423_ _07970_ _07936_ vssd1 vssd1 vccd1 vccd1 _08125_ sky130_fd_sc_hd__or4_1
X_12723_ _05292_ _05299_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__xor2_1
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16491_ _09099_ _09100_ vssd1 vssd1 vccd1 vccd1 _09101_ sky130_fd_sc_hd__or2_1
XFILLER_203_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18230_ rbzero.wall_tracer.trackDistY\[-11\] _01996_ _02007_ _09286_ vssd1 vssd1
+ vccd1 vccd1 _00566_ sky130_fd_sc_hd__o22a_1
X_15442_ _08053_ _08055_ vssd1 vssd1 vccd1 vccd1 _08056_ sky130_fd_sc_hd__xnor2_1
X_12654_ _05218_ _05342_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__xnor2_2
XFILLER_43_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11605_ _04319_ _04320_ _04321_ _03932_ _03946_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__o221a_1
X_18161_ _07827_ _07914_ _01876_ _01940_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__o31a_1
XFILLER_145_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15373_ _07508_ _07542_ _07549_ _07593_ vssd1 vssd1 vccd1 vccd1 _07987_ sky130_fd_sc_hd__or4_1
XFILLER_169_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12585_ rbzero.wall_tracer.visualWallDist\[2\] _03815_ vssd1 vssd1 vccd1 vccd1 _05274_
+ sky130_fd_sc_hd__nor2_1
XFILLER_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17112_ _09527_ _09565_ _09563_ vssd1 vssd1 vccd1 vccd1 _09652_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14324_ _06789_ _06793_ _06965_ vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__o21ba_1
X_11536_ rbzero.debug_overlay.vplaneX\[-4\] _04242_ _04209_ rbzero.debug_overlay.vplaneX\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__a22o_1
X_18092_ _01737_ _01738_ _01740_ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__a21bo_1
XFILLER_102_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17043_ _09582_ _09583_ vssd1 vssd1 vccd1 vccd1 _09584_ sky130_fd_sc_hd__and2b_1
X_14255_ _06933_ _06939_ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__nand2_1
XFILLER_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11467_ _04183_ _04184_ _03910_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__mux2_1
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ _05618_ _05745_ _05635_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__a21o_1
XFILLER_87_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10418_ _03421_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14186_ _06853_ _06873_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__nor2_1
XFILLER_178_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11398_ _03826_ _04109_ _04115_ _04116_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__a211o_1
XFILLER_180_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13137_ _05809_ _05811_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__and2b_1
XFILLER_135_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ rbzero.tex_r1\[50\] rbzero.tex_r1\[51\] _03377_ vssd1 vssd1 vccd1 vccd1 _03385_
+ sky130_fd_sc_hd__mux2_1
X_18994_ _02657_ vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17945_ _01721_ _01727_ rbzero.wall_tracer.trackDistX\[8\] _09276_ vssd1 vssd1 vccd1
+ vccd1 _00561_ sky130_fd_sc_hd__o2bb2a_1
X_13068_ _05742_ _05755_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__and2_1
XFILLER_112_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12019_ net8 _04727_ _04718_ net5 vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__and4bb_1
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17876_ _01657_ _01658_ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__nand2_1
XFILLER_152_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19615_ _02753_ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__buf_4
XFILLER_226_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16827_ _09096_ _09098_ _09234_ _09368_ vssd1 vssd1 vccd1 vccd1 _09369_ sky130_fd_sc_hd__o31ai_4
XFILLER_113_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19546_ rbzero.pov.spi_buffer\[68\] rbzero.pov.spi_buffer\[69\] _02932_ vssd1 vssd1
+ vccd1 vccd1 _02942_ sky130_fd_sc_hd__mux2_1
XFILLER_207_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16758_ _09303_ _09307_ _09308_ _09283_ vssd1 vssd1 vccd1 vccd1 _09309_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15709_ _08286_ _08309_ vssd1 vssd1 vccd1 vccd1 _08323_ sky130_fd_sc_hd__xnor2_1
X_19477_ rbzero.pov.spi_buffer\[35\] rbzero.pov.spi_buffer\[36\] _02899_ vssd1 vssd1
+ vccd1 vccd1 _02906_ sky130_fd_sc_hd__mux2_1
XFILLER_55_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16689_ rbzero.traced_texa\[-7\] _09262_ _09263_ rbzero.wall_tracer.visualWallDist\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__a22o_1
XFILLER_224_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18428_ rbzero.wall_tracer.rayAddendX\[-3\] _02179_ _03812_ vssd1 vssd1 vccd1 vccd1
+ _02180_ sky130_fd_sc_hd__mux2_1
XFILLER_210_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18359_ _04999_ _02001_ _02118_ vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__a21oi_1
XFILLER_187_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21370_ _00393_ _01386_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20321_ rbzero.traced_texVinit\[10\] _03260_ _09267_ _09764_ vssd1 vssd1 vccd1 vccd1
+ _01404_ sky130_fd_sc_hd__a22o_1
XFILLER_200_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20252_ _03254_ vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__clkinv_2
XFILLER_66_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20183_ _03200_ _03203_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__nand2_1
XFILLER_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12370_ _05061_ _05062_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__nand2_1
XFILLER_138_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11321_ _04038_ _03919_ _03953_ _04039_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__or4_1
X_20519_ net129 _00535_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14040_ _06710_ _06728_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__xnor2_1
XFILLER_180_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11252_ rbzero.tex_r0\[41\] _03964_ _03965_ _03932_ vssd1 vssd1 vccd1 vccd1 _03971_
+ sky130_fd_sc_hd__a31o_1
XFILLER_84_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10203_ _03308_ vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11183_ _03859_ _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__nand2_1
XTAP_6421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ _07742_ _07800_ _08603_ vssd1 vssd1 vccd1 vccd1 _08604_ sky130_fd_sc_hd__o21ai_1
XTAP_5720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17730_ _01496_ _10152_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__or2b_1
XTAP_6487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14942_ _07551_ _07555_ vssd1 vssd1 vccd1 vccd1 _07556_ sky130_fd_sc_hd__nand2_1
XFILLER_121_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17661_ _10163_ _10164_ _01444_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__nand3_1
XTAP_5797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14873_ _07378_ _07387_ _07399_ _07423_ vssd1 vssd1 vccd1 vccd1 _07487_ sky130_fd_sc_hd__or4_1
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19400_ _02864_ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__clkbuf_4
X_16612_ _09075_ _09077_ vssd1 vssd1 vccd1 vccd1 _09221_ sky130_fd_sc_hd__and2_1
XFILLER_169_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13824_ _06471_ _06472_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__nand2_1
XFILLER_91_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17592_ _10126_ _10127_ _10109_ vssd1 vssd1 vccd1 vccd1 _10129_ sky130_fd_sc_hd__a21oi_1
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19331_ _02856_ vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__clkinv_2
XFILLER_56_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16543_ _09149_ _09151_ vssd1 vssd1 vccd1 vccd1 _09152_ sky130_fd_sc_hd__nor2_1
XFILLER_245_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13755_ _06442_ _06438_ vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__or2b_1
X_10967_ _03711_ vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12706_ _05255_ _05384_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__xnor2_1
X_19262_ _02815_ vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16474_ _09081_ _09082_ _09013_ vssd1 vssd1 vccd1 vccd1 _09084_ sky130_fd_sc_hd__a21o_1
XFILLER_149_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13686_ _06309_ _06327_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__nand2_1
X_10898_ _03675_ vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__clkbuf_1
X_18213_ _01991_ _01992_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__xnor2_1
X_15425_ _07443_ _07708_ vssd1 vssd1 vccd1 vccd1 _08039_ sky130_fd_sc_hd__nor2_1
XFILLER_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12637_ _05204_ _05271_ _05305_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__o21ai_1
X_19193_ rbzero.spi_registers.new_vshift\[0\] _02775_ vssd1 vssd1 vccd1 vccd1 _02776_
+ sky130_fd_sc_hd__or2_1
XFILLER_180_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18144_ _01906_ _01907_ _01904_ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__o21a_1
XFILLER_191_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15356_ _04928_ _07698_ vssd1 vssd1 vccd1 vccd1 _07970_ sky130_fd_sc_hd__nand2_2
X_12568_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__or2_1
XFILLER_106_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14307_ _06571_ _06973_ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__xor2_1
XFILLER_129_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11519_ _03783_ _04223_ _04207_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__and3_2
X_18075_ _01736_ _01751_ _01855_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__a21bo_1
XFILLER_144_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15287_ _07876_ _07877_ _07899_ vssd1 vssd1 vccd1 vccd1 _07901_ sky130_fd_sc_hd__nand3_1
X_12499_ _03816_ _05069_ _05112_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__nand3_2
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17026_ _09438_ _09440_ vssd1 vssd1 vccd1 vccd1 _09567_ sky130_fd_sc_hd__nor2_1
X_14238_ _06911_ _06926_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__or2_1
XFILLER_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14169_ _05660_ _06482_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__or2_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _02648_ vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17928_ _01708_ _01710_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__or2_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17859_ _01640_ _01641_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__xor2_1
XFILLER_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20870_ net54 _00886_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19529_ _02933_ vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_241_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21353_ _00376_ _01369_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20304_ _03258_ vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__clkinv_2
XFILLER_107_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21284_ _00333_ _01300_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_100_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20235_ rbzero.traced_texa\[11\] rbzero.texV\[11\] vssd1 vssd1 vccd1 vccd1 _03250_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_116_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20166_ _03093_ _03191_ _03192_ _03064_ rbzero.texV\[-1\] vssd1 vssd1 vccd1 vccd1
+ _01317_ sky130_fd_sc_hd__a32o_1
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20097_ rbzero.traced_texa\[-12\] rbzero.texV\[-12\] vssd1 vssd1 vccd1 vccd1 _03135_
+ sky130_fd_sc_hd__nand2_1
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _04581_ _04582_ _04583_ _03909_ _03944_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__o221a_1
XFILLER_217_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ rbzero.tex_g0\[21\] rbzero.tex_g0\[20\] _03627_ vssd1 vssd1 vccd1 vccd1 _03635_
+ sky130_fd_sc_hd__mux2_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20999_ net55 _01015_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13540_ _06193_ _06208_ _06191_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__a21bo_1
X_10752_ _03598_ vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13471_ _05979_ _06025_ _06159_ _05980_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__a211oi_1
XFILLER_158_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10683_ _03562_ vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15210_ _07818_ _07823_ _07519_ vssd1 vssd1 vccd1 vccd1 _07824_ sky130_fd_sc_hd__a21o_2
XFILLER_185_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12422_ rbzero.map_rom.c6 _05114_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__and2_1
XFILLER_16_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16190_ _08792_ _08801_ vssd1 vssd1 vccd1 vccd1 _08802_ sky130_fd_sc_hd__xnor2_1
XFILLER_205_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15141_ _07746_ _07754_ vssd1 vssd1 vccd1 vccd1 _07755_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12353_ rbzero.debug_overlay.facingY\[-5\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__or2_1
XFILLER_51_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11304_ rbzero.tex_r0\[1\] rbzero.tex_r0\[0\] _03936_ vssd1 vssd1 vccd1 vccd1 _04023_
+ sky130_fd_sc_hd__mux2_1
X_15072_ _07453_ rbzero.wall_tracer.stepDistY\[4\] vssd1 vssd1 vccd1 vccd1 _07686_
+ sky130_fd_sc_hd__and2_1
XFILLER_154_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12284_ _04977_ rbzero.wall_tracer.trackDistY\[-6\] vssd1 vssd1 vccd1 vccd1 _04978_
+ sky130_fd_sc_hd__nor2_1
XFILLER_177_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14023_ _06703_ _06711_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__and2_1
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18900_ _02607_ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__clkbuf_4
XFILLER_84_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11235_ _03953_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__buf_4
X_19880_ _03110_ vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__clkinv_2
XFILLER_49_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18831_ _02428_ _02535_ _02549_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__a21o_1
XTAP_6240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11166_ rbzero.traced_texVinit\[9\] rbzero.texV\[9\] _03880_ _03881_ vssd1 vssd1
+ vccd1 vccd1 _03885_ sky130_fd_sc_hd__a22o_1
XTAP_6251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18762_ _02166_ _02484_ _02485_ _02158_ rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__a32o_1
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15974_ rbzero.wall_tracer.texu\[0\] _07338_ _07266_ _08587_ vssd1 vssd1 vccd1 vccd1
+ _00481_ sky130_fd_sc_hd__o211a_1
X_11097_ rbzero.wall_tracer.state\[0\] vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__inv_2
XTAP_5561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17713_ _10150_ _10151_ _01497_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__a21o_2
XTAP_5572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14925_ _07492_ _07538_ vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__nand2_1
XTAP_5594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18693_ _02416_ _02417_ _02418_ _02407_ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__a22o_1
XFILLER_236_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17644_ _01427_ _01428_ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__and2_1
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14856_ _07435_ vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__clkbuf_4
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13807_ _06458_ _06477_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__xor2_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17575_ _08771_ _09611_ _09732_ _08046_ vssd1 vssd1 vccd1 vccd1 _10112_ sky130_fd_sc_hd__a22o_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14787_ _07388_ _07400_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__nor2_1
XFILLER_51_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11999_ net42 _04694_ _04697_ net44 vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__a22o_1
XFILLER_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19314_ _02846_ _02847_ vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__nor2_1
X_16526_ _09133_ _09134_ vssd1 vssd1 vccd1 vccd1 _09135_ sky130_fd_sc_hd__or2_1
XFILLER_225_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13738_ _06425_ _06426_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19245_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.new_leak\[1\] _02804_
+ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__mux2_1
X_16457_ _08935_ _08933_ vssd1 vssd1 vccd1 vccd1 _09067_ sky130_fd_sc_hd__and2b_1
XFILLER_176_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13669_ _06323_ _06335_ _06356_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__or3_1
XFILLER_73_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15408_ _08019_ _08020_ _08021_ vssd1 vssd1 vccd1 vccd1 _08022_ sky130_fd_sc_hd__a21boi_1
XFILLER_121_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19176_ _09247_ _02764_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__and2_1
X_16388_ _08274_ _07621_ _08671_ _08592_ vssd1 vssd1 vccd1 vccd1 _08998_ sky130_fd_sc_hd__o22a_1
XFILLER_157_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18127_ _01906_ _01907_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15339_ _07932_ _07950_ vssd1 vssd1 vccd1 vccd1 _07953_ sky130_fd_sc_hd__nor2_1
XFILLER_145_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18058_ _09163_ _09611_ _01837_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__a21oi_1
XFILLER_201_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17009_ _09548_ _09549_ vssd1 vssd1 vccd1 vccd1 _09550_ sky130_fd_sc_hd__nand2_1
XFILLER_132_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20020_ _03124_ vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__clkinv_2
XFILLER_99_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20922_ net74 _00938_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20853_ _00071_ _00869_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20784_ net102 _00800_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21405_ net114 _01421_ vssd1 vssd1 vccd1 vccd1 gpout3.clk_div\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21336_ _00359_ _01352_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21267_ _00316_ _01283_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_235_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11020_ rbzero.map_rom.b6 rbzero.map_rom.a6 rbzero.map_rom.i_row\[4\] vssd1 vssd1
+ vccd1 vccd1 _03748_ sky130_fd_sc_hd__or3_1
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20218_ _03234_ _03235_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__and2b_1
XFILLER_132_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21198_ _00247_ _01214_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20149_ rbzero.traced_texa\[-3\] rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1 _03178_
+ sky130_fd_sc_hd__nand2_1
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _05659_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__clkbuf_4
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _07329_ vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__clkbuf_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _03288_ _04592_ _04631_ _04632_ net9 _04625_ vssd1 vssd1 vccd1 vccd1 _04633_
+ sky130_fd_sc_hd__mux4_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15690_ _08292_ _08299_ vssd1 vssd1 vccd1 vccd1 _08304_ sky130_fd_sc_hd__and2b_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14641_ _05001_ _07254_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__nor2_1
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11853_ _03909_ _04564_ _04565_ _04566_ _03919_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__o221a_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17360_ _09895_ _09896_ _09897_ vssd1 vssd1 vccd1 vccd1 _09898_ sky130_fd_sc_hd__nor3_1
X_10804_ rbzero.tex_g0\[29\] rbzero.tex_g0\[28\] _03616_ vssd1 vssd1 vccd1 vccd1 _03626_
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14572_ _06991_ _07006_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__nand2_1
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11784_ rbzero.tex_b0\[2\] _03959_ _03916_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__a21o_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16311_ _08918_ _08921_ _04938_ vssd1 vssd1 vccd1 vccd1 _08922_ sky130_fd_sc_hd__a21o_1
XFILLER_198_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13523_ _05858_ _05868_ _06211_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__a21oi_1
X_17291_ _08594_ _08595_ _09829_ _08628_ vssd1 vssd1 vccd1 vccd1 _09830_ sky130_fd_sc_hd__or4_1
XFILLER_186_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10735_ _03589_ vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19030_ _02676_ vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16242_ _07625_ _08852_ vssd1 vssd1 vccd1 vccd1 _08853_ sky130_fd_sc_hd__or2_1
XFILLER_174_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13454_ _06114_ _06120_ _06098_ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__o21ai_1
X_10666_ rbzero.tex_g1\[30\] rbzero.tex_g1\[31\] _03552_ vssd1 vssd1 vccd1 vccd1 _03554_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12405_ rbzero.wall_tracer.rayAddendY\[-4\] _05091_ _05093_ _05097_ vssd1 vssd1 vccd1
+ vccd1 _05098_ sky130_fd_sc_hd__or4_1
XFILLER_51_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16173_ _08781_ _08784_ _07519_ vssd1 vssd1 vccd1 vccd1 _08785_ sky130_fd_sc_hd__a21o_1
X_13385_ _05699_ _05738_ _06071_ _06072_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__a22o_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10597_ _03517_ vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15124_ _07728_ _07737_ vssd1 vssd1 vccd1 vccd1 _07738_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12336_ _05029_ vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12267_ rbzero.wall_tracer.trackDistX\[3\] _04941_ _04943_ _04960_ vssd1 vssd1 vccd1
+ vccd1 _04961_ sky130_fd_sc_hd__a22o_1
X_15055_ _07342_ _05267_ _07668_ _04932_ vssd1 vssd1 vccd1 vccd1 _07669_ sky130_fd_sc_hd__a211o_1
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19932_ _03116_ vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__clkinv_2
XFILLER_218_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14006_ _06650_ _06653_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__xor2_1
X_11218_ rbzero.tex_r0\[58\] _03936_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__and2_1
XFILLER_214_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19863_ _03109_ vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__clkinv_2
XFILLER_218_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12198_ net43 _04899_ _04900_ net44 vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__a22o_1
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11149_ _03846_ _03864_ _03867_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__o21a_1
X_18814_ _02524_ _02525_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__or2b_1
XTAP_6070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19794_ _04104_ _03094_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__and2_1
XTAP_6081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18745_ _02458_ _02459_ _02468_ _02469_ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__o22ai_1
XTAP_5380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15957_ _08568_ _08570_ vssd1 vssd1 vccd1 vccd1 _08571_ sky130_fd_sc_hd__xnor2_4
XFILLER_114_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14908_ _07501_ _07508_ _07520_ _07521_ vssd1 vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18676_ rbzero.wall_tracer.rayAddendY\[-3\] _02405_ _03812_ vssd1 vssd1 vccd1 vccd1
+ _02406_ sky130_fd_sc_hd__mux2_1
XFILLER_97_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15888_ _08498_ _08499_ _08500_ vssd1 vssd1 vccd1 vccd1 _08502_ sky130_fd_sc_hd__a21o_1
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17627_ _10107_ _10093_ vssd1 vssd1 vccd1 vccd1 _10163_ sky130_fd_sc_hd__or2b_1
XFILLER_224_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14839_ _07351_ vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__buf_4
XFILLER_149_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17558_ _07840_ vssd1 vssd1 vccd1 vccd1 _10095_ sky130_fd_sc_hd__clkbuf_4
XFILLER_205_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16509_ _09010_ _09109_ _09117_ vssd1 vssd1 vccd1 vccd1 _09118_ sky130_fd_sc_hd__a21oi_1
XFILLER_204_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17489_ _04940_ _10026_ vssd1 vssd1 vccd1 vccd1 _10027_ sky130_fd_sc_hd__nand2_1
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19228_ _02796_ vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__clkbuf_1
XFILLER_177_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19159_ rbzero.spi_registers.new_sky\[0\] rbzero.spi_registers.got_new_sky _02724_
+ _02753_ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__a31o_1
XFILLER_145_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21121_ _00170_ _01137_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_236_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21052_ _00101_ _01068_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_232_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20003_ _03114_ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__buf_4
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20905_ net67 _00921_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[42\] sky130_fd_sc_hd__dfxtp_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20836_ _00054_ _00852_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20767_ net100 _00783_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10520_ rbzero.tex_r0\[36\] rbzero.tex_r0\[35\] _03468_ vssd1 vssd1 vccd1 vccd1 _03477_
+ sky130_fd_sc_hd__mux2_1
XFILLER_211_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20698_ net101 _00714_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_183_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10451_ rbzero.tex_r1\[2\] rbzero.tex_r1\[3\] _03433_ vssd1 vssd1 vccd1 vccd1 _03439_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13170_ _05553_ _05722_ _05768_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__and3_1
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10382_ rbzero.tex_r1\[35\] rbzero.tex_r1\[36\] _03400_ vssd1 vssd1 vccd1 vccd1 _03403_
+ sky130_fd_sc_hd__mux2_1
XFILLER_164_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12121_ _04820_ o_rgb[23] _04827_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__a21bo_1
XFILLER_87_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21319_ _00342_ _01335_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12052_ net42 _04750_ _04755_ net44 vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a22o_1
XFILLER_111_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11003_ rbzero.wall_tracer.state\[1\] vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__inv_2
X_16860_ _09391_ _09400_ vssd1 vssd1 vccd1 vccd1 _09402_ sky130_fd_sc_hd__or2_1
XFILLER_215_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15811_ _08422_ _08423_ vssd1 vssd1 vccd1 vccd1 _08425_ sky130_fd_sc_hd__xnor2_1
XFILLER_237_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16791_ rbzero.wall_tracer.trackDistX\[-5\] _09301_ _09331_ _09337_ vssd1 vssd1 vccd1
+ vccd1 _00548_ sky130_fd_sc_hd__o22a_1
XFILLER_111_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18530_ _02247_ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__buf_2
XFILLER_234_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15742_ _08330_ _08348_ vssd1 vssd1 vccd1 vccd1 _08356_ sky130_fd_sc_hd__xor2_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _05621_ _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__nor2_1
XFILLER_133_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _04611_ _04519_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__nor2_1
X_18461_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.debug_overlay.vplaneX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__nor2_1
XFILLER_94_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15673_ _08263_ _08265_ vssd1 vssd1 vccd1 vccd1 _08287_ sky130_fd_sc_hd__xnor2_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _05501_ _05571_ _05573_ _05405_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__o211a_1
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17412_ _09913_ _09949_ vssd1 vssd1 vccd1 vccd1 _09950_ sky130_fd_sc_hd__xnor2_1
XFILLER_221_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _04950_ _07246_ _07249_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__o21ai_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ rbzero.tex_b1\[34\] _03934_ _03928_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__a21o_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18392_ rbzero.debug_overlay.vplaneX\[-7\] rbzero.wall_tracer.rayAddendX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__nor2_1
XFILLER_92_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _09776_ _09881_ vssd1 vssd1 vccd1 vccd1 _09882_ sky130_fd_sc_hd__xor2_1
XFILLER_53_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14555_ rbzero.wall_tracer.stepDistY\[6\] _07225_ _07193_ vssd1 vssd1 vccd1 vccd1
+ _07226_ sky130_fd_sc_hd__mux2_1
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ rbzero.tex_b0\[27\] rbzero.tex_b0\[26\] _04013_ vssd1 vssd1 vccd1 vccd1 _04482_
+ sky130_fd_sc_hd__mux2_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13506_ _05739_ _05852_ _06194_ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__a21bo_1
X_17274_ _09166_ _08735_ vssd1 vssd1 vccd1 vccd1 _09813_ sky130_fd_sc_hd__nor2_1
X_10718_ rbzero.tex_g1\[5\] rbzero.tex_g1\[6\] _03574_ vssd1 vssd1 vccd1 vccd1 _03581_
+ sky130_fd_sc_hd__mux2_1
XFILLER_187_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14486_ _05447_ _07169_ _05602_ vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__a21o_1
XFILLER_158_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11698_ rbzero.tex_g1\[58\] _04374_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__and2_1
X_19013_ _02667_ vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__clkbuf_1
X_16225_ _07338_ _08836_ vssd1 vssd1 vccd1 vccd1 _08837_ sky130_fd_sc_hd__nand2_1
XFILLER_228_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13437_ _06124_ _06125_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__xnor2_1
X_10649_ rbzero.tex_g1\[38\] rbzero.tex_g1\[39\] _03541_ vssd1 vssd1 vccd1 vccd1 _03545_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16156_ _08619_ _08618_ vssd1 vssd1 vccd1 vccd1 _08768_ sky130_fd_sc_hd__nand2_1
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13368_ _06038_ _06056_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15107_ _07472_ _07664_ vssd1 vssd1 vccd1 vccd1 _07721_ sky130_fd_sc_hd__nor2_1
XFILLER_177_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12319_ _05000_ _05012_ _04993_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__o21a_1
XFILLER_170_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16087_ _08588_ _08699_ vssd1 vssd1 vccd1 vccd1 _08700_ sky130_fd_sc_hd__xnor2_4
X_13299_ _05941_ _05985_ _05986_ _05987_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__a22o_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15038_ _07260_ _07351_ vssd1 vssd1 vccd1 vccd1 _07652_ sky130_fd_sc_hd__nor2_2
XFILLER_130_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19915_ _03114_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__buf_4
XFILLER_170_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19846_ _03107_ vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__clkinv_2
XFILLER_190_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16989_ _08510_ _08850_ vssd1 vssd1 vccd1 vccd1 _09530_ sky130_fd_sc_hd__nor2_1
X_19777_ _03083_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__inv_2
XFILLER_68_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18728_ rbzero.wall_tracer.rayAddendY\[1\] _02197_ _02453_ _02157_ vssd1 vssd1 vccd1
+ vccd1 _02454_ sky130_fd_sc_hd__a22o_1
XFILLER_209_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18659_ _02386_ _02387_ _02389_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__or3_1
XFILLER_97_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20621_ net79 _00637_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20552_ net120 _00568_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20483_ net111 _00499_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21104_ _00153_ _01120_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_6817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout100 net104 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__buf_2
Xfanout111 net113 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_2
XFILLER_248_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout122 net126 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__buf_2
XFILLER_248_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout133 net134 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_2
X_21035_ _00084_ _01051_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_232_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12670_ _05310_ _05322_ _05353_ _05358_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__and4_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ rbzero.tex_g0\[51\] rbzero.tex_g0\[50\] _03935_ vssd1 vssd1 vccd1 vccd1 _04338_
+ sky130_fd_sc_hd__mux2_1
X_20819_ _00037_ _00835_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14340_ _05458_ vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__buf_2
X_11552_ rbzero.debug_overlay.facingY\[-2\] _04245_ _04243_ rbzero.debug_overlay.facingY\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__a22o_1
XFILLER_195_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10503_ _03445_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__clkbuf_4
X_14271_ _06877_ _06879_ _06840_ vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__a21oi_1
XFILLER_155_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11483_ _03780_ _04200_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__nand2_1
XFILLER_109_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16010_ _08616_ _08622_ vssd1 vssd1 vccd1 vccd1 _08623_ sky130_fd_sc_hd__xor2_1
X_13222_ _05591_ _05672_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__or2_1
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10434_ rbzero.tex_r1\[10\] rbzero.tex_r1\[11\] _03422_ vssd1 vssd1 vccd1 vccd1 _03430_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13153_ _05840_ _05841_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__nand2_1
X_10365_ rbzero.tex_r1\[43\] rbzero.tex_r1\[44\] _03389_ vssd1 vssd1 vccd1 vccd1 _03394_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12104_ net51 _04798_ _04799_ net53 _04811_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__a221o_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17961_ _08240_ _08241_ _09976_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__a21oi_1
X_13084_ _05729_ _05772_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _03357_ vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16912_ _09452_ _09453_ vssd1 vssd1 vccd1 vccd1 _09454_ sky130_fd_sc_hd__nand2_1
XFILLER_215_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19700_ _02728_ _03054_ vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__nand2_1
X_12035_ net6 net7 _04743_ net8 vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a22oi_1
X_17892_ _09955_ _07914_ _01673_ vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__o21ai_1
XFILLER_214_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16843_ _07878_ _08850_ vssd1 vssd1 vccd1 vccd1 _09385_ sky130_fd_sc_hd__nor2_1
X_19631_ rbzero.pov.ready_buffer\[72\] _02963_ _03001_ vssd1 vssd1 vccd1 vccd1 _03002_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_226_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19562_ rbzero.pov.ss_buffer\[1\] rbzero.pov.ss_buffer\[0\] _09243_ vssd1 vssd1 vccd1
+ vccd1 _02950_ sky130_fd_sc_hd__mux2_1
X_16774_ _09303_ _09321_ _09322_ _09282_ vssd1 vssd1 vccd1 vccd1 _09323_ sky130_fd_sc_hd__a31o_1
XFILLER_111_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13986_ _06662_ _06674_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18513_ _02248_ _02250_ _02257_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__a21oi_1
X_15725_ _08333_ _08334_ _08338_ vssd1 vssd1 vccd1 vccd1 _08339_ sky130_fd_sc_hd__a21o_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12937_ _05489_ _05612_ _05625_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__a21o_1
X_19493_ _02914_ vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18444_ _02181_ _02190_ _02192_ _02193_ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__and4_1
XFILLER_221_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15656_ _08245_ _08269_ vssd1 vssd1 vccd1 vccd1 _08270_ sky130_fd_sc_hd__xor2_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12868_ _05499_ _05521_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__nor2_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14607_ rbzero.wall_tracer.trackDistX\[-7\] rbzero.wall_tracer.trackDistY\[-7\] _07258_
+ vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__mux2_1
X_18375_ rbzero.wall_tracer.trackDistY\[10\] rbzero.wall_tracer.stepDistY\[10\] vssd1
+ vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__xnor2_1
X_11819_ _03908_ _04530_ _04531_ _04532_ _03944_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__o221a_1
X_15587_ _08199_ _08200_ vssd1 vssd1 vccd1 vccd1 _08201_ sky130_fd_sc_hd__xor2_2
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12799_ _05447_ _05479_ _05482_ _05487_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__o22a_2
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17326_ _09863_ _09864_ vssd1 vssd1 vccd1 vccd1 _09865_ sky130_fd_sc_hd__and2b_1
X_14538_ rbzero.wall_tracer.stepDistY\[3\] _07211_ _07193_ vssd1 vssd1 vccd1 vccd1
+ _07212_ sky130_fd_sc_hd__mux2_1
XFILLER_159_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17257_ _09794_ _09795_ vssd1 vssd1 vccd1 vccd1 _09796_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14469_ _05577_ _07150_ _07154_ _05602_ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__a211oi_1
XFILLER_175_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16208_ _08684_ _08659_ vssd1 vssd1 vccd1 vccd1 _08820_ sky130_fd_sc_hd__or2b_1
XFILLER_174_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17188_ _08779_ _09611_ vssd1 vssd1 vccd1 vccd1 _09728_ sky130_fd_sc_hd__nand2_1
XFILLER_143_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16139_ _07469_ _08067_ _07520_ _08750_ vssd1 vssd1 vccd1 vccd1 _08751_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_196_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19829_ _03106_ vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__clkinv_2
XFILLER_233_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20604_ net81 _00620_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_205_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20535_ net131 _00551_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20466_ net119 _00482_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20397_ net138 _00428_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21018_ net80 _01034_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_done sky130_fd_sc_hd__dfxtp_2
XTAP_5957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13840_ _06527_ _06528_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13771_ _06408_ _06459_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__xor2_1
XFILLER_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10983_ rbzero.tex_b0\[8\] rbzero.tex_b0\[7\] _03715_ vssd1 vssd1 vccd1 vccd1 _03720_
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15510_ _07435_ _07423_ _08123_ _07698_ vssd1 vssd1 vccd1 vccd1 _08124_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12722_ _05402_ _05323_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__nand2_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16490_ rbzero.debug_overlay.playerY\[-2\] rbzero.debug_overlay.playerX\[-2\] _07343_
+ vssd1 vssd1 vccd1 vccd1 _09100_ sky130_fd_sc_hd__mux2_1
XFILLER_188_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15441_ _07997_ _08054_ vssd1 vssd1 vccd1 vccd1 _08055_ sky130_fd_sc_hd__and2_1
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12653_ _05338_ _05339_ _05340_ _05341_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__a31o_1
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18160_ _01874_ _01875_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__nand2_1
XFILLER_180_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11604_ rbzero.tex_g0\[1\] rbzero.tex_g0\[0\] _03936_ vssd1 vssd1 vccd1 vccd1 _04321_
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15372_ _07985_ vssd1 vssd1 vccd1 vccd1 _07986_ sky130_fd_sc_hd__buf_2
XFILLER_180_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12584_ _05182_ _05272_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__xnor2_2
XFILLER_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17111_ _09376_ _09525_ _09523_ vssd1 vssd1 vccd1 vccd1 _09651_ sky130_fd_sc_hd__a21o_1
X_14323_ _06788_ _06841_ _07008_ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__a21oi_1
X_18091_ _01782_ _01783_ _01785_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__a21bo_1
XFILLER_141_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11535_ rbzero.debug_overlay.vplaneX\[-5\] _04214_ _04237_ rbzero.debug_overlay.vplaneX\[-6\]
+ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__a22o_1
XFILLER_184_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17042_ _09580_ _09581_ vssd1 vssd1 vccd1 vccd1 _09583_ sky130_fd_sc_hd__nand2_1
XFILLER_221_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14254_ _06940_ _06942_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__nor2_1
XFILLER_176_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11466_ rbzero.tex_r1\[7\] rbzero.tex_r1\[6\] _04168_ vssd1 vssd1 vccd1 vccd1 _04184_
+ sky130_fd_sc_hd__mux2_1
XFILLER_109_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13205_ _05629_ _05609_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__or2_1
X_10417_ rbzero.tex_r1\[18\] rbzero.tex_r1\[19\] _03411_ vssd1 vssd1 vccd1 vccd1 _03421_
+ sky130_fd_sc_hd__mux2_1
X_14185_ _06853_ _06873_ vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__and2_1
X_11397_ _03291_ _03294_ _03295_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__o21a_2
XFILLER_125_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13136_ _05822_ _05824_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__or2b_1
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _03384_ vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_225_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18993_ rbzero.pov.spi_buffer\[44\] rbzero.pov.ready_buffer\[44\] _02651_ vssd1 vssd1
+ vccd1 vccd1 _02657_ sky130_fd_sc_hd__mux2_1
XFILLER_112_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17944_ _09279_ _01726_ _09283_ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__a21oi_1
X_13067_ _05742_ _05755_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__nor2_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _03348_ vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_238_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12018_ _04717_ _04519_ _04726_ net6 net7 vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__o2111a_1
XFILLER_66_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17875_ _07678_ _08531_ _01535_ vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__o21ai_1
XFILLER_61_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19614_ rbzero.pov.ready_buffer\[69\] _02963_ _02981_ _02987_ vssd1 vssd1 vccd1 vccd1
+ _02988_ sky130_fd_sc_hd__o211a_1
XFILLER_66_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16826_ _09235_ _09233_ _09232_ vssd1 vssd1 vccd1 vccd1 _09368_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16757_ _09304_ _09305_ _09306_ vssd1 vssd1 vccd1 vccd1 _09308_ sky130_fd_sc_hd__a21o_1
X_19545_ _02941_ vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13969_ _06639_ _06657_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15708_ _08221_ _08321_ vssd1 vssd1 vccd1 vccd1 _08322_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16688_ rbzero.traced_texa\[-8\] _09262_ _09263_ rbzero.wall_tracer.visualWallDist\[-8\]
+ vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__a22o_1
X_19476_ _02905_ vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15639_ _07571_ _07572_ _07573_ _07645_ vssd1 vssd1 vccd1 vccd1 _08253_ sky130_fd_sc_hd__a211o_1
XFILLER_146_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18427_ _09256_ _02170_ _02171_ _02178_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__a31o_1
XFILLER_94_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18358_ _02116_ _02117_ _01612_ _01995_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__o211a_1
XFILLER_159_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17309_ _09846_ _09847_ vssd1 vssd1 vccd1 vccd1 _09848_ sky130_fd_sc_hd__and2_1
XFILLER_187_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18289_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.stepDistY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__nor2_1
XFILLER_124_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20320_ rbzero.traced_texVinit\[9\] _03260_ _09267_ _09640_ vssd1 vssd1 vccd1 vccd1
+ _01403_ sky130_fd_sc_hd__a22o_1
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20251_ _03254_ vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__clkinv_2
XFILLER_196_1280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20182_ rbzero.traced_texa\[2\] rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1 _03206_
+ sky130_fd_sc_hd__nand2_1
XFILLER_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11320_ _04026_ _03908_ _03898_ _04030_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__or4_1
X_20518_ net132 _00534_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11251_ rbzero.tex_r0\[40\] _03962_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__and2_1
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20449_ net118 _00000_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10202_ rbzero.tex_b1\[56\] rbzero.tex_b1\[57\] _03300_ vssd1 vssd1 vccd1 vccd1 _03308_
+ sky130_fd_sc_hd__mux2_1
XTAP_7134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11182_ _03855_ _03858_ _03893_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__a21oi_2
XTAP_7145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15990_ _07552_ _07736_ vssd1 vssd1 vccd1 vccd1 _08603_ sky130_fd_sc_hd__or2_1
XTAP_5710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14941_ _07424_ _07552_ _07553_ _07554_ vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17660_ _10163_ _10164_ _01444_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__a21o_1
XTAP_5787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14872_ _07416_ _07485_ vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__nor2_1
XFILLER_76_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16611_ _09181_ _09219_ vssd1 vssd1 vccd1 vccd1 _09220_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13823_ _06440_ _06510_ _06511_ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__o21a_1
XFILLER_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17591_ _10109_ _10126_ _10127_ vssd1 vssd1 vccd1 vccd1 _10128_ sky130_fd_sc_hd__and3_1
XFILLER_1_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16542_ _08995_ _09002_ _09150_ vssd1 vssd1 vccd1 vccd1 _09151_ sky130_fd_sc_hd__a21oi_1
X_19330_ _02856_ vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__clkinv_2
X_13754_ _06438_ _06442_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__xnor2_1
XFILLER_182_1302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10966_ rbzero.tex_b0\[16\] rbzero.tex_b0\[15\] _03704_ vssd1 vssd1 vccd1 vccd1 _03711_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ _05253_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__inv_2
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19261_ rbzero.spi_registers.new_other\[1\] rbzero.spi_registers.spi_buffer\[1\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__mux2_1
X_16473_ _09013_ _09081_ _09082_ vssd1 vssd1 vccd1 vccd1 _09083_ sky130_fd_sc_hd__nand3_1
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13685_ _06329_ _06373_ _05434_ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__a21oi_1
X_10897_ rbzero.tex_b0\[49\] rbzero.tex_b0\[48\] _03671_ vssd1 vssd1 vccd1 vccd1 _03675_
+ sky130_fd_sc_hd__mux2_1
XFILLER_245_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18212_ rbzero.wall_tracer.trackDistX\[11\] rbzero.wall_tracer.stepDistX\[11\] vssd1
+ vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__xor2_1
X_15424_ _07435_ _07387_ vssd1 vssd1 vccd1 vccd1 _08038_ sky130_fd_sc_hd__or2_1
XFILLER_148_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12636_ _05199_ _05324_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__xor2_4
X_19192_ rbzero.spi_registers.got_new_vshift _02724_ vssd1 vssd1 vccd1 vccd1 _02775_
+ sky130_fd_sc_hd__nand2_1
XFILLER_223_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18143_ _01856_ _01886_ _01922_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__a21bo_1
XFILLER_157_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15355_ _07435_ _07355_ vssd1 vssd1 vccd1 vccd1 _07969_ sky130_fd_sc_hd__or2_1
X_12567_ _05251_ _05253_ _05255_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__or3_1
XFILLER_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14306_ _05432_ _06992_ _06994_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__a21o_1
XFILLER_141_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18074_ _01752_ _01735_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__or2b_1
X_11518_ _04230_ _04231_ _04234_ _04235_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__or4_2
X_15286_ _07876_ _07877_ _07899_ vssd1 vssd1 vccd1 vccd1 _07900_ sky130_fd_sc_hd__a21o_1
XFILLER_141_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12498_ _03790_ _05186_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__nand2_1
X_17025_ _09527_ _09565_ vssd1 vssd1 vccd1 vccd1 _09566_ sky130_fd_sc_hd__xor2_1
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14237_ _06913_ _06919_ _06925_ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__o21a_1
X_11449_ _04165_ _04166_ _03916_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__mux2_1
XFILLER_125_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14168_ _06820_ _06856_ vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__nand2_1
XFILLER_152_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _05803_ _05806_ _05807_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__a21bo_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _06786_ _06787_ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__nor2_1
X_18976_ rbzero.pov.spi_buffer\[36\] rbzero.pov.ready_buffer\[36\] _02640_ vssd1 vssd1
+ vccd1 vccd1 _02648_ sky130_fd_sc_hd__mux2_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _01603_ _01604_ _01709_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__o21a_1
XFILLER_113_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17858_ _01575_ _01577_ _01458_ _01574_ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_187_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16809_ _04947_ _09283_ _09353_ vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__a21oi_1
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17789_ _01571_ _01572_ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__and2_1
XFILLER_241_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19528_ rbzero.pov.spi_buffer\[59\] rbzero.pov.spi_buffer\[60\] _02932_ vssd1 vssd1
+ vccd1 vccd1 _02933_ sky130_fd_sc_hd__mux2_1
XFILLER_207_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19459_ _02896_ vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21352_ _00375_ _01368_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20303_ _03258_ vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__clkinv_2
XFILLER_198_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21283_ _00332_ _01299_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20234_ _09245_ _03248_ _03249_ _03064_ rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1
+ _01328_ sky130_fd_sc_hd__a32o_1
XFILLER_122_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20165_ _03188_ _03189_ _03183_ _03187_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__a211o_1
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20096_ _03134_ vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _03634_ vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20998_ net59 _01014_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10751_ rbzero.tex_g0\[54\] rbzero.tex_g0\[53\] _03593_ vssd1 vssd1 vccd1 vccd1 _03598_
+ sky130_fd_sc_hd__mux2_1
XFILLER_242_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13470_ _05978_ _05979_ _06025_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__nor3_1
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10682_ rbzero.tex_g1\[22\] rbzero.tex_g1\[23\] _03552_ vssd1 vssd1 vccd1 vccd1 _03562_
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12421_ _05113_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__buf_4
XFILLER_142_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15140_ _07747_ _07753_ vssd1 vssd1 vccd1 vccd1 _07754_ sky130_fd_sc_hd__xor2_1
XFILLER_166_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12352_ rbzero.debug_overlay.facingY\[-5\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__nand2_1
XFILLER_166_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11303_ rbzero.tex_r0\[2\] _04001_ _03942_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__a21o_1
X_15071_ _07684_ vssd1 vssd1 vccd1 vccd1 _07685_ sky130_fd_sc_hd__buf_2
X_12283_ rbzero.wall_tracer.trackDistX\[-6\] vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__inv_2
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14022_ _06697_ _06702_ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__nand2_1
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11234_ _03872_ _03894_ _03952_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__nor3_2
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18830_ _02547_ _02548_ _02535_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__a21oi_1
XTAP_6230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11165_ _03876_ _03877_ _03882_ _03883_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__o22ai_1
XTAP_6241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15973_ _07338_ _08586_ vssd1 vssd1 vccd1 vccd1 _08587_ sky130_fd_sc_hd__nand2_1
X_11096_ _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__clkbuf_4
XFILLER_122_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18761_ _02482_ _02483_ _02461_ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__o21ai_1
XTAP_6285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17712_ _10152_ _01496_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__xor2_1
XTAP_5573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14924_ rbzero.debug_overlay.playerX\[-3\] _07411_ vssd1 vssd1 vccd1 vccd1 _07538_
+ sky130_fd_sc_hd__nand2_1
XFILLER_23_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18692_ _02419_ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__inv_2
XTAP_5595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17643_ _10169_ _01426_ vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__or2_1
X_14855_ _07355_ vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__buf_2
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13806_ _06489_ _06494_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__xnor2_1
X_17574_ _08779_ _09857_ _09465_ vssd1 vssd1 vccd1 vccd1 _10111_ sky130_fd_sc_hd__a21bo_4
X_14786_ _07399_ vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__buf_4
XFILLER_56_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11998_ _04664_ net15 _04116_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__and3_1
XFILLER_189_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16525_ _07515_ _08723_ _08986_ _08987_ vssd1 vssd1 vccd1 vccd1 _09134_ sky130_fd_sc_hd__o31a_1
X_19313_ rbzero.pov.spi_counter\[2\] _02840_ _02838_ vssd1 vssd1 vccd1 vccd1 _02847_
+ sky130_fd_sc_hd__o21ai_1
X_13737_ _06317_ _06388_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__nor2_1
XFILLER_108_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10949_ rbzero.tex_b0\[24\] rbzero.tex_b0\[23\] _03693_ vssd1 vssd1 vccd1 vccd1 _03702_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16456_ _09063_ _09064_ _09054_ vssd1 vssd1 vccd1 vccd1 _09066_ sky130_fd_sc_hd__a21o_1
XFILLER_143_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19244_ _02805_ vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__clkbuf_1
X_13668_ _06323_ _06356_ _06335_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__o21ai_1
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15407_ _07945_ _08006_ _08018_ vssd1 vssd1 vccd1 vccd1 _08021_ sky130_fd_sc_hd__nand3_1
XFILLER_160_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12619_ rbzero.wall_tracer.visualWallDist\[10\] _03816_ _03790_ rbzero.wall_tracer.visualWallDist\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__or4b_1
X_19175_ rbzero.spi_registers.new_floor\[0\] rbzero.color_floor\[0\] _02763_ vssd1
+ vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__mux2_1
X_16387_ _08599_ _07916_ vssd1 vssd1 vccd1 vccd1 _08997_ sky130_fd_sc_hd__nor2_1
X_13599_ _06262_ _06287_ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__xnor2_4
XFILLER_247_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18126_ _01695_ _01810_ _01808_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__a21oi_1
XFILLER_160_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15338_ _07614_ _07590_ vssd1 vssd1 vccd1 vccd1 _07952_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18057_ _09163_ _09611_ _01837_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__and3_1
X_15269_ _07554_ _07793_ _07520_ _07882_ vssd1 vssd1 vccd1 vccd1 _07883_ sky130_fd_sc_hd__a22o_1
XFILLER_144_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17008_ _07620_ _09166_ _08536_ _09018_ vssd1 vssd1 vccd1 vccd1 _09549_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_160_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18959_ rbzero.pov.spi_buffer\[28\] rbzero.pov.ready_buffer\[28\] _02629_ vssd1 vssd1
+ vccd1 vccd1 _02639_ sky130_fd_sc_hd__mux2_1
XFILLER_79_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20921_ net68 _00937_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20852_ _00070_ _00868_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20783_ net102 _00799_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_other
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21404_ net114 _01420_ vssd1 vssd1 vccd1 vccd1 gpout3.clk_div\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21335_ _00358_ _01351_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21266_ _00315_ _01282_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20217_ rbzero.traced_texa\[8\] rbzero.texV\[8\] vssd1 vssd1 vccd1 vccd1 _03235_
+ sky130_fd_sc_hd__nand2_1
X_21197_ _00246_ _01213_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20148_ rbzero.traced_texa\[-3\] rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1 _03177_
+ sky130_fd_sc_hd__or2_1
XFILLER_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12970_ _05489_ _05628_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__xnor2_1
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20079_ _03130_ vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__clkinv_2
XFILLER_218_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ gpout0.vpos\[1\] vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__buf_2
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ rbzero.wall_tracer.visualWallDist\[3\] _07253_ _07288_ _07289_ _07266_ vssd1
+ vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__o221a_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ rbzero.tex_b1\[31\] _03938_ _03940_ _03928_ vssd1 vssd1 vccd1 vccd1 _04566_
+ sky130_fd_sc_hd__a31o_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _03625_ vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__clkbuf_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14571_ _07238_ vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ rbzero.tex_b0\[3\] _04143_ _04145_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__and3_1
XFILLER_57_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16310_ _07338_ _08919_ _08920_ _07694_ vssd1 vssd1 vccd1 vccd1 _08921_ sky130_fd_sc_hd__o31ai_4
XFILLER_198_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13522_ _05775_ _05869_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__nor2_1
XFILLER_242_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17290_ _04933_ _07648_ _07650_ vssd1 vssd1 vccd1 vccd1 _09829_ sky130_fd_sc_hd__a21oi_4
XFILLER_159_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10734_ rbzero.tex_g0\[62\] rbzero.tex_g0\[61\] _03512_ vssd1 vssd1 vccd1 vccd1 _03589_
+ sky130_fd_sc_hd__mux2_1
XFILLER_207_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16241_ _08851_ vssd1 vssd1 vccd1 vccd1 _08852_ sky130_fd_sc_hd__clkbuf_4
X_13453_ _06123_ _06135_ _06140_ _06141_ vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__a31o_1
XFILLER_16_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10665_ _03553_ vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12404_ rbzero.wall_tracer.rayAddendY\[-3\] rbzero.wall_tracer.rayAddendY\[-2\] _05095_
+ _05096_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__or4_1
X_16172_ _04933_ _08782_ _08783_ _07822_ vssd1 vssd1 vccd1 vccd1 _08784_ sky130_fd_sc_hd__a31o_1
XFILLER_142_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13384_ _05699_ _05738_ _06071_ _06072_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__nand4_2
XFILLER_142_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10596_ rbzero.tex_g1\[63\] net49 _03433_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__mux2_1
XFILLER_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15123_ _07468_ _07736_ vssd1 vssd1 vccd1 vccd1 _07737_ sky130_fd_sc_hd__nor2_1
XFILLER_86_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12335_ _04934_ rbzero.map_rom.d6 _05028_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__mux2_1
XFILLER_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15054_ _07341_ _05110_ vssd1 vssd1 vccd1 vccd1 _07668_ sky130_fd_sc_hd__nor2_1
XFILLER_147_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19931_ _03116_ vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__clkinv_2
XFILLER_177_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12266_ _04946_ _04958_ _04959_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__a21o_1
XFILLER_108_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14005_ _06407_ _06691_ _06692_ _06693_ vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__a22o_1
X_11217_ _03935_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__buf_4
X_19862_ _03109_ vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__clkinv_2
X_12197_ net49 net40 net39 net41 net34 _04874_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__mux4_1
XFILLER_214_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18813_ _02530_ _02531_ _02528_ _02529_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__o211ai_1
XTAP_6060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11148_ _03866_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__inv_2
XTAP_6071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19793_ _03094_ _03095_ vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__nor2_1
XFILLER_233_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18744_ _02465_ _02467_ _09256_ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__o21ai_1
XTAP_5370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15956_ _08110_ _08569_ vssd1 vssd1 vccd1 vccd1 _08570_ sky130_fd_sc_hd__and2_1
X_11079_ _03290_ gpout0.hpos\[8\] gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _03802_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_37_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14907_ _07352_ _07512_ _07515_ vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__or3b_4
X_15887_ _08498_ _08499_ _08500_ vssd1 vssd1 vccd1 vccd1 _08501_ sky130_fd_sc_hd__nand3_1
XFILLER_23_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18675_ _09256_ _02396_ _02397_ _02404_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a31o_1
XFILLER_237_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17626_ _10070_ _10085_ _10083_ vssd1 vssd1 vccd1 vccd1 _10162_ sky130_fd_sc_hd__a21o_1
X_14838_ _07342_ _05080_ vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__or2_1
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17557_ _08594_ _08595_ _07840_ _08917_ vssd1 vssd1 vccd1 vccd1 _10094_ sky130_fd_sc_hd__or4_1
X_14769_ _07341_ _05230_ _07382_ _04932_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__a211o_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16508_ _09112_ _09116_ vssd1 vssd1 vccd1 vccd1 _09117_ sky130_fd_sc_hd__xnor2_1
XFILLER_204_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17488_ _10020_ _10025_ vssd1 vssd1 vccd1 vccd1 _10026_ sky130_fd_sc_hd__or2_1
XFILLER_225_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19227_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.new_floor\[0\]
+ _02795_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__mux2_1
X_16439_ _07229_ _07234_ _07237_ _08474_ _07241_ vssd1 vssd1 vccd1 vccd1 _09049_ sky130_fd_sc_hd__o41a_1
XFILLER_34_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19158_ _03442_ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__buf_4
XFILLER_195_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18109_ _01754_ _01755_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__nor2_1
XFILLER_173_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19089_ _03442_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__buf_6
XFILLER_172_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21120_ _00169_ _01136_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21051_ _00100_ _01067_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20002_ _03122_ vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__clkinv_2
XFILLER_236_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20904_ net67 _00920_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20835_ _00053_ _00851_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_243_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20766_ net100 _00782_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20697_ net101 _00713_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_195_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10450_ _03438_ vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10381_ _03402_ vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12120_ _04820_ _04519_ net31 net30 vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__o211a_1
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21318_ _00341_ _01334_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12051_ o_tex_oeb0 _04755_ _04759_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__a21o_1
X_21249_ _00298_ _01265_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_215_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11002_ _03729_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__buf_4
XFILLER_46_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15810_ _08422_ _08423_ vssd1 vssd1 vccd1 vccd1 _08424_ sky130_fd_sc_hd__nand2_1
XFILLER_63_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16790_ _09303_ _09335_ _09336_ _09282_ vssd1 vssd1 vccd1 vccd1 _09337_ sky130_fd_sc_hd__a31o_1
XFILLER_120_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15741_ _08353_ _08354_ vssd1 vssd1 vccd1 vccd1 _08355_ sky130_fd_sc_hd__nand2_1
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12953_ _05641_ _05632_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__nand2_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11904_ net12 net13 vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__nand2_1
XFILLER_233_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15672_ _08283_ _08285_ vssd1 vssd1 vccd1 vccd1 _08286_ sky130_fd_sc_hd__nor2_1
X_18460_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.debug_overlay.vplaneX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__and2_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12884_ _05357_ _05430_ _05572_ _05462_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__a211o_1
XFILLER_2_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _09947_ _09948_ vssd1 vssd1 vccd1 vccd1 _09949_ sky130_fd_sc_hd__nand2_1
X_14623_ _04954_ _07254_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__nor2_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11835_ rbzero.tex_b1\[35\] _03859_ _03901_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__and3_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18391_ _02143_ _02144_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__and2b_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _09878_ _09880_ vssd1 vssd1 vccd1 vccd1 _09881_ sky130_fd_sc_hd__xnor2_1
XFILLER_202_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14554_ _07223_ _07096_ _07213_ _07224_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__o211ai_2
XFILLER_187_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _03954_ _04455_ _04463_ _04480_ _03896_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__a311o_1
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13505_ _05853_ _05846_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__or2b_1
XFILLER_159_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17273_ _09810_ _09811_ vssd1 vssd1 vccd1 vccd1 _09812_ sky130_fd_sc_hd__nand2_1
X_10717_ _03580_ vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__clkbuf_1
X_14485_ _07130_ _07030_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__nand2_1
XFILLER_174_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11697_ rbzero.tex_g1\[57\] rbzero.tex_g1\[56\] _04378_ vssd1 vssd1 vccd1 vccd1 _04413_
+ sky130_fd_sc_hd__mux2_1
XFILLER_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16224_ _08585_ _08835_ vssd1 vssd1 vccd1 vccd1 _08836_ sky130_fd_sc_hd__xnor2_1
X_19012_ rbzero.pov.spi_buffer\[53\] rbzero.pov.ready_buffer\[53\] _02662_ vssd1 vssd1
+ vccd1 vccd1 _02667_ sky130_fd_sc_hd__mux2_1
XFILLER_186_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13436_ _06112_ _06111_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__or2b_1
XFILLER_31_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10648_ _03544_ vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16155_ _08747_ _08766_ vssd1 vssd1 vccd1 vccd1 _08767_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13367_ _06040_ _06054_ _06055_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__o21a_1
X_10579_ rbzero.tex_r0\[8\] rbzero.tex_r0\[7\] _03501_ vssd1 vssd1 vccd1 vccd1 _03508_
+ sky130_fd_sc_hd__mux2_1
XFILLER_154_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15106_ _07717_ _07719_ vssd1 vssd1 vccd1 vccd1 _07720_ sky130_fd_sc_hd__xor2_1
X_12318_ _05003_ _05007_ _05005_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__o21a_1
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16086_ _08697_ _08698_ vssd1 vssd1 vccd1 vccd1 _08699_ sky130_fd_sc_hd__nand2_2
XFILLER_181_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13298_ _05941_ _05985_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__xor2_1
XFILLER_108_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15037_ _04933_ _07648_ _07650_ vssd1 vssd1 vccd1 vccd1 _07651_ sky130_fd_sc_hd__a21o_4
X_19914_ _04702_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__buf_4
X_12249_ rbzero.wall_tracer.trackDistX\[3\] _04941_ rbzero.wall_tracer.trackDistX\[2\]
+ _04942_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__o22a_1
XFILLER_29_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19845_ _03107_ vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__clkinv_2
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19776_ gpout0.vpos\[8\] gpout0.vpos\[7\] _03076_ _03082_ vssd1 vssd1 vccd1 vccd1
+ _03083_ sky130_fd_sc_hd__or4_1
XFILLER_111_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16988_ _07878_ _08978_ vssd1 vssd1 vccd1 vccd1 _09529_ sky130_fd_sc_hd__or2_1
X_18727_ _02436_ _02452_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__xnor2_1
X_15939_ _08529_ _08552_ vssd1 vssd1 vccd1 vccd1 _08553_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18658_ _02371_ _02382_ _02388_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__o21ai_1
XFILLER_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17609_ _10035_ _10026_ _10145_ vssd1 vssd1 vccd1 vccd1 _10146_ sky130_fd_sc_hd__and3_1
XFILLER_184_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18589_ _02327_ _02328_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__and2_1
XFILLER_212_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20620_ net79 _00636_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20551_ net120 _00567_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20482_ net111 _00498_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21103_ _00152_ _01119_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_6818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout101 net104 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__buf_2
XFILLER_99_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout112 net113 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__buf_2
Xfanout123 net124 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__buf_2
X_21034_ _00083_ _01050_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[2\] sky130_fd_sc_hd__dfxtp_1
Xfanout134 net140 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_2
XFILLER_102_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ rbzero.tex_g0\[49\] rbzero.tex_g0\[48\] _04148_ vssd1 vssd1 vccd1 vccd1 _04337_
+ sky130_fd_sc_hd__mux2_1
XFILLER_179_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20818_ _00036_ _00834_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11551_ rbzero.debug_overlay.facingY\[-4\] _04242_ _04209_ rbzero.debug_overlay.facingY\[-3\]
+ _04268_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__a221o_1
XFILLER_180_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20749_ net104 _00765_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10502_ _03467_ vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__clkbuf_1
X_14270_ _06879_ _06880_ _06956_ _06958_ vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__and4_2
X_11482_ _04196_ _04199_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__nor2_1
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13221_ _05795_ _05797_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10433_ _03429_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13152_ _05783_ _05781_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__or2b_1
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10364_ _03393_ vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12103_ net52 _04773_ _04768_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__and3_1
XFILLER_124_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17960_ _01740_ _01741_ vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__and2_1
X_13083_ _05616_ _05726_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__nor2_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10295_ rbzero.tex_b1\[12\] rbzero.tex_b1\[13\] _03355_ vssd1 vssd1 vccd1 vccd1 _03357_
+ sky130_fd_sc_hd__mux2_1
XFILLER_219_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16911_ _09449_ _08917_ _09188_ vssd1 vssd1 vccd1 vccd1 _09453_ sky130_fd_sc_hd__o21ai_1
X_12034_ net5 _04735_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__nor2_1
XFILLER_78_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17891_ _09955_ _07914_ _01673_ vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__or3_1
XFILLER_120_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19630_ _02833_ _03000_ _02981_ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__o21a_1
X_16842_ _09177_ _09162_ vssd1 vssd1 vccd1 vccd1 _09384_ sky130_fd_sc_hd__and2b_1
XFILLER_215_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19561_ _02949_ vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__clkbuf_1
X_13985_ _06664_ _06672_ _06673_ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__a21bo_1
X_16773_ _09318_ _09319_ _09320_ vssd1 vssd1 vccd1 vccd1 _09322_ sky130_fd_sc_hd__a21o_1
XFILLER_65_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18512_ _02247_ rbzero.wall_tracer.rayAddendX\[4\] vssd1 vssd1 vccd1 vccd1 _02257_
+ sky130_fd_sc_hd__xnor2_1
X_15724_ _07879_ _07843_ _08336_ _08337_ vssd1 vssd1 vccd1 vccd1 _08338_ sky130_fd_sc_hd__o31ai_1
X_12936_ _05470_ _05514_ _05520_ _05447_ _05524_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__a221o_4
XFILLER_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19492_ rbzero.pov.spi_buffer\[42\] rbzero.pov.spi_buffer\[43\] _02910_ vssd1 vssd1
+ vccd1 vccd1 _02914_ sky130_fd_sc_hd__mux2_1
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18443_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] _02184_
+ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__a21o_1
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15655_ _08247_ _08267_ _08268_ vssd1 vssd1 vccd1 vccd1 _08269_ sky130_fd_sc_hd__a21boi_1
X_12867_ _05497_ _05554_ _05555_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__a21o_1
XFILLER_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14606_ rbzero.wall_tracer.visualWallDist\[-8\] _07253_ _07264_ _07265_ _07266_ vssd1
+ vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__o221a_1
X_11818_ rbzero.tex_b1\[59\] _03859_ _03901_ _03914_ vssd1 vssd1 vccd1 vccd1 _04532_
+ sky130_fd_sc_hd__a31o_1
XFILLER_221_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18374_ _02125_ _02127_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__nand2_1
X_15586_ _07260_ _07408_ _07356_ _07420_ vssd1 vssd1 vccd1 vccd1 _08200_ sky130_fd_sc_hd__or4_2
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12798_ _05483_ _05486_ _05460_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__mux2_2
XFILLER_159_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _09859_ _09860_ _09862_ vssd1 vssd1 vccd1 vccd1 _09864_ sky130_fd_sc_hd__a21o_1
XFILLER_226_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14537_ _07100_ _07210_ vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__nand2_1
XFILLER_239_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11749_ rbzero.tex_b0\[45\] rbzero.tex_b0\[44\] _03980_ vssd1 vssd1 vccd1 vccd1 _04464_
+ sky130_fd_sc_hd__mux2_1
XFILLER_105_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17256_ _07882_ _09115_ vssd1 vssd1 vccd1 vccd1 _09795_ sky130_fd_sc_hd__nor2_1
X_14468_ _05527_ _07151_ _07153_ _05535_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__o211a_1
XFILLER_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16207_ _08817_ _08818_ vssd1 vssd1 vccd1 vccd1 _08819_ sky130_fd_sc_hd__nand2_1
X_13419_ _05625_ _05959_ _06107_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__or3b_1
X_17187_ _09718_ _09726_ vssd1 vssd1 vccd1 vccd1 _09727_ sky130_fd_sc_hd__xor2_1
X_14399_ _05531_ _07055_ _07087_ vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__o21ai_1
XFILLER_143_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16138_ _07384_ _07385_ vssd1 vssd1 vccd1 vccd1 _08750_ sky130_fd_sc_hd__nand2_2
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16069_ _08680_ _08681_ vssd1 vssd1 vccd1 vccd1 _08682_ sky130_fd_sc_hd__xor2_1
XFILLER_115_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19828_ _03106_ vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__clkinv_2
XFILLER_57_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19759_ rbzero.pov.ready_buffer\[9\] _03060_ _03062_ _02428_ _03015_ vssd1 vssd1
+ vccd1 vccd1 _01032_ sky130_fd_sc_hd__a221o_1
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20603_ net81 _00619_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20534_ net130 _00550_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20465_ net128 _00481_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20396_ net138 _00427_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21017_ net81 _01033_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_212_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13770_ _06412_ _06413_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__xnor2_1
X_10982_ _03719_ vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12721_ _05356_ _05397_ _05409_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__nand3b_2
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15440_ _07994_ _07996_ vssd1 vssd1 vccd1 vccd1 _08054_ sky130_fd_sc_hd__or2_1
X_12652_ _05220_ _05294_ _05280_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__a21oi_2
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11603_ rbzero.tex_g0\[2\] _04013_ _04014_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__a21o_1
X_15371_ _07529_ _07984_ vssd1 vssd1 vccd1 vccd1 _07985_ sky130_fd_sc_hd__and2_1
XFILLER_141_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12583_ _05179_ _05181_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__nand2_1
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17110_ _09634_ _09516_ vssd1 vssd1 vccd1 vccd1 _09650_ sky130_fd_sc_hd__or2b_1
X_14322_ _05431_ _07010_ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__nor2_1
XFILLER_180_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18090_ _01861_ _01870_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__xnor2_1
X_11534_ _04104_ _04102_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__nor2_2
XFILLER_129_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17041_ _09580_ _09581_ vssd1 vssd1 vccd1 vccd1 _09582_ sky130_fd_sc_hd__nor2_1
XFILLER_184_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14253_ _06930_ _06941_ vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__nand2_1
XFILLER_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11465_ rbzero.tex_r1\[5\] rbzero.tex_r1\[4\] _04168_ vssd1 vssd1 vccd1 vccd1 _04183_
+ sky130_fd_sc_hd__mux2_1
XFILLER_184_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13204_ _05618_ _05745_ _05625_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__a21o_1
XFILLER_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10416_ _03420_ vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__clkbuf_1
X_14184_ _06855_ _06872_ _06870_ vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__a21oi_1
XFILLER_178_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11396_ _04111_ _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__nand2_4
X_13135_ _05823_ _05709_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10347_ rbzero.tex_r1\[51\] rbzero.tex_r1\[52\] _03377_ vssd1 vssd1 vccd1 vccd1 _03384_
+ sky130_fd_sc_hd__mux2_1
X_18992_ _02656_ vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__clkbuf_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _01724_ _01725_ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__xnor2_1
X_13066_ _05743_ _05754_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10278_ rbzero.tex_b1\[20\] rbzero.tex_b1\[21\] _03344_ vssd1 vssd1 vccd1 vccd1 _03348_
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12017_ _04717_ o_rgb[23] vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__nand2_1
XFILLER_6_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17874_ _07678_ _08531_ _01535_ vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__or3_1
XFILLER_152_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19613_ rbzero.debug_overlay.playerX\[1\] _02982_ _02986_ vssd1 vssd1 vccd1 vccd1
+ _02987_ sky130_fd_sc_hd__a21o_1
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16825_ _09361_ _09367_ rbzero.wall_tracer.trackDistX\[-1\] _09276_ vssd1 vssd1 vccd1
+ vccd1 _00552_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_241_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19544_ rbzero.pov.spi_buffer\[67\] rbzero.pov.spi_buffer\[68\] _02932_ vssd1 vssd1
+ vccd1 vccd1 _02941_ sky130_fd_sc_hd__mux2_1
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16756_ _09304_ _09305_ _09306_ vssd1 vssd1 vccd1 vccd1 _09307_ sky130_fd_sc_hd__nand3_1
XFILLER_47_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13968_ _06641_ _06656_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__xor2_1
XFILLER_111_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15707_ _08320_ _08319_ vssd1 vssd1 vccd1 vccd1 _08321_ sky130_fd_sc_hd__nor2_1
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12919_ _05591_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__clkbuf_4
X_19475_ rbzero.pov.spi_buffer\[34\] rbzero.pov.spi_buffer\[35\] _02899_ vssd1 vssd1
+ vccd1 vccd1 _02905_ sky130_fd_sc_hd__mux2_1
XFILLER_222_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13899_ _06435_ _06331_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__nor2_1
X_16687_ rbzero.traced_texa\[-9\] _09262_ _09263_ rbzero.wall_tracer.visualWallDist\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18426_ _09256_ _02177_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__nor2_1
X_15638_ _08201_ _08203_ vssd1 vssd1 vccd1 vccd1 _08252_ sky130_fd_sc_hd__xnor2_2
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18357_ _02113_ _02114_ _02115_ _04940_ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__a31o_1
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15569_ _08180_ _08181_ _08182_ vssd1 vssd1 vccd1 vccd1 _08183_ sky130_fd_sc_hd__a21bo_1
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17308_ _09826_ _09845_ vssd1 vssd1 vccd1 vccd1 _09847_ sky130_fd_sc_hd__or2_1
XFILLER_174_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18288_ _07275_ _02001_ _02057_ vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__a21oi_1
XFILLER_148_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17239_ _09696_ _09661_ vssd1 vssd1 vccd1 vccd1 _09778_ sky130_fd_sc_hd__or2b_1
XFILLER_190_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20250_ _03125_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__buf_4
XFILLER_127_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20181_ rbzero.traced_texa\[2\] rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1 _03205_
+ sky130_fd_sc_hd__or2_1
XFILLER_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20517_ net132 _00533_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11250_ rbzero.tex_r0\[43\] rbzero.tex_r0\[42\] _03959_ vssd1 vssd1 vccd1 vccd1 _03969_
+ sky130_fd_sc_hd__mux2_1
X_20448_ net123 _00015_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10201_ _03307_ vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__clkbuf_1
XTAP_7124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11181_ _03899_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__buf_4
XFILLER_49_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20379_ net116 _00410_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14940_ _07481_ _07482_ _07483_ vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__a21oi_4
XTAP_6489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14871_ _07484_ vssd1 vssd1 vccd1 vccd1 _07485_ sky130_fd_sc_hd__buf_2
XTAP_5799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16610_ _09217_ _09218_ vssd1 vssd1 vccd1 vccd1 _09219_ sky130_fd_sc_hd__xor2_1
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13822_ _05641_ _06305_ _06321_ _05738_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__a22o_1
X_17590_ _10122_ _10123_ _10125_ vssd1 vssd1 vccd1 vccd1 _10127_ sky130_fd_sc_hd__a21o_1
XFILLER_112_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16541_ _08886_ _08889_ _09001_ vssd1 vssd1 vccd1 vccd1 _09150_ sky130_fd_sc_hd__a21oi_1
X_13753_ _06439_ _06441_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__or2b_1
XFILLER_21_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10965_ _03710_ vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12704_ _05361_ _05363_ _05382_ _05392_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__o31a_1
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19260_ _02814_ vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__clkbuf_1
XFILLER_245_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16472_ _09077_ _09078_ _09080_ vssd1 vssd1 vccd1 vccd1 _09082_ sky130_fd_sc_hd__a21o_1
XFILLER_189_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13684_ _06309_ _06315_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__nand2_1
XFILLER_95_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10896_ _03674_ vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18211_ rbzero.wall_tracer.trackDistX\[10\] rbzero.wall_tracer.stepDistX\[10\] _01919_
+ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__a21o_1
XFILLER_54_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15423_ _07467_ _07423_ vssd1 vssd1 vccd1 vccd1 _08037_ sky130_fd_sc_hd__nor2_1
X_12635_ _05204_ _05271_ _05276_ _05296_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__o31a_1
X_19191_ _02773_ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__clkbuf_2
XFILLER_54_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18142_ _01887_ _01854_ vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__or2b_1
XFILLER_169_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15354_ _07965_ _07966_ _07967_ vssd1 vssd1 vccd1 vccd1 _07968_ sky130_fd_sc_hd__a21o_1
XFILLER_157_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12566_ rbzero.wall_tracer.rayAddendX\[-3\] _05254_ _05219_ vssd1 vssd1 vccd1 vccd1
+ _05255_ sky130_fd_sc_hd__mux2_2
XFILLER_196_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14305_ _06981_ _06993_ vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__and2_1
X_11517_ _04223_ _04233_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__and2_1
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18073_ _01779_ _01794_ _01792_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__a21o_1
X_15285_ _07888_ _07898_ vssd1 vssd1 vccd1 vccd1 _07899_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12497_ _05143_ _05184_ _05185_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__a21oi_4
X_17024_ _09563_ _09564_ vssd1 vssd1 vccd1 vccd1 _09565_ sky130_fd_sc_hd__nor2_1
X_14236_ _06923_ _06924_ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__nand2_1
X_11448_ rbzero.tex_r1\[25\] rbzero.tex_r1\[24\] _03904_ vssd1 vssd1 vccd1 vccd1 _04166_
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14167_ _05668_ _06222_ _06341_ _06819_ vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__a31o_1
XFILLER_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11379_ _04040_ _04097_ rbzero.row_render.vinf vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13118_ _05715_ _05804_ _05749_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__or3_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _06785_ _06783_ _06784_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__and3_1
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18975_ _02647_ vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__clkbuf_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17926_ _01605_ _01515_ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__or2b_1
X_13049_ _05634_ _05636_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__nand2_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17857_ _01638_ _01639_ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16808_ _09345_ _09349_ _09350_ _09275_ _09352_ vssd1 vssd1 vccd1 vccd1 _09353_ sky130_fd_sc_hd__o311a_1
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17788_ _07631_ _07827_ _01570_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__o21ai_1
XFILLER_208_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19527_ _02864_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__clkbuf_4
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16739_ rbzero.wall_tracer.trackDistX\[-11\] _09276_ _09286_ _09291_ vssd1 vssd1
+ vccd1 vccd1 _00542_ sky130_fd_sc_hd__o22a_1
XFILLER_35_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19458_ rbzero.pov.spi_buffer\[26\] rbzero.pov.spi_buffer\[27\] _02888_ vssd1 vssd1
+ vccd1 vccd1 _02896_ sky130_fd_sc_hd__mux2_1
XFILLER_195_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18409_ _02143_ _02155_ _02144_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__o21ai_1
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19389_ _02861_ vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__clkinv_2
XFILLER_188_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21351_ _00374_ _01367_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20302_ _03258_ vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__clkinv_2
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21282_ _00331_ _01298_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20233_ _03240_ _03245_ _03246_ _03247_ vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__nand4_1
XFILLER_157_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20164_ _03190_ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__inv_2
XFILLER_130_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20095_ _09247_ _03132_ _03133_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__and3_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20997_ net56 _01013_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_168_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ _03597_ vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10681_ _03561_ vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_205_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12420_ _05073_ _05111_ _05112_ _05069_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_139_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12351_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__or2_1
XFILLER_103_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ rbzero.tex_r0\[3\] _03939_ _03941_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__and3_1
X_15070_ _07672_ _07673_ vssd1 vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__and2_1
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12282_ _04962_ rbzero.wall_tracer.trackDistY\[-7\] vssd1 vssd1 vccd1 vccd1 _04976_
+ sky130_fd_sc_hd__nor2_1
XFILLER_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14021_ _06661_ _06675_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11233_ _03871_ _03840_ _03868_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__nor3_1
XFILLER_181_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11164_ rbzero.texV\[8\] _03875_ _03873_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__a21oi_1
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18760_ _02461_ _02482_ _02483_ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__or3_1
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15972_ _08583_ _08585_ vssd1 vssd1 vccd1 vccd1 _08586_ sky130_fd_sc_hd__xnor2_1
X_11095_ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__buf_2
XTAP_6286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17711_ _01494_ _01495_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__xnor2_1
XTAP_6297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14923_ rbzero.debug_overlay.playerX\[-3\] vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__inv_2
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18691_ _02407_ _02416_ _02417_ _02418_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__and4_1
XTAP_5585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17642_ _10169_ _01426_ vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__nand2_1
X_14854_ _07467_ vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__clkbuf_4
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13805_ _06491_ _06493_ vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__xor2_1
XFILLER_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17573_ _09979_ _09981_ vssd1 vssd1 vccd1 vccd1 _10110_ sky130_fd_sc_hd__nand2_1
XFILLER_189_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14785_ _07398_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__clkbuf_4
XFILLER_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11997_ o_tex_oeb0 _04697_ _04698_ net47 _04706_ vssd1 vssd1 vccd1 vccd1 _04707_
+ sky130_fd_sc_hd__a221o_1
XFILLER_216_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19312_ rbzero.pov.spi_counter\[2\] _02840_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__and2_1
XFILLER_72_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16524_ _09129_ _09132_ vssd1 vssd1 vccd1 vccd1 _09133_ sky130_fd_sc_hd__xnor2_1
XFILLER_205_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13736_ _05767_ _06343_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__nor2_1
XFILLER_188_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10948_ _03701_ vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19243_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.new_leak\[0\] _02804_
+ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__mux2_1
X_16455_ _09054_ _09063_ _09064_ vssd1 vssd1 vccd1 vccd1 _09065_ sky130_fd_sc_hd__nand3_1
XFILLER_188_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13667_ _06316_ _06322_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__nor2_1
XFILLER_143_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10879_ _03665_ vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15406_ _07968_ _07978_ vssd1 vssd1 vccd1 vccd1 _08020_ sky130_fd_sc_hd__xor2_1
X_12618_ _05303_ _05306_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__xnor2_1
X_19174_ rbzero.spi_registers.got_new_floor _02720_ vssd1 vssd1 vccd1 vccd1 _02763_
+ sky130_fd_sc_hd__nand2_2
X_16386_ _08886_ _08889_ vssd1 vssd1 vccd1 vccd1 _08996_ sky130_fd_sc_hd__nand2_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13598_ _06285_ _06286_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__nor2_2
XFILLER_160_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18125_ _01904_ _01905_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__nand2_1
XFILLER_247_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15337_ _07932_ _07950_ vssd1 vssd1 vccd1 vccd1 _07951_ sky130_fd_sc_hd__xor2_1
X_12549_ rbzero.wall_tracer.visualWallDist\[-6\] _05189_ rbzero.wall_tracer.rcp_sel\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__a21o_1
XFILLER_121_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18056_ _09428_ _08923_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__nor2_1
XANTENNA_1 _01823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15268_ _07571_ _07572_ vssd1 vssd1 vccd1 vccd1 _07882_ sky130_fd_sc_hd__nand2_2
XFILLER_172_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17007_ _08086_ _07620_ _07936_ _08671_ vssd1 vssd1 vccd1 vccd1 _09548_ sky130_fd_sc_hd__or4_1
X_14219_ _06901_ _06907_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__nand2_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15199_ _07783_ _07812_ vssd1 vssd1 vccd1 vccd1 _07813_ sky130_fd_sc_hd__and2_1
XFILLER_125_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18958_ _02638_ vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17909_ _01563_ _01525_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__or2b_1
X_18889_ rbzero.spi_registers.spi_counter\[4\] _02597_ vssd1 vssd1 vccd1 vccd1 _02600_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_41_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20920_ net67 _00936_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20851_ _00069_ _00867_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20782_ net88 _00798_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21403_ net106 _01419_ vssd1 vssd1 vccd1 vccd1 gpout2.clk_div\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21334_ _00357_ _01350_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21265_ _00314_ _01281_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_237_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20216_ rbzero.traced_texa\[8\] rbzero.texV\[8\] vssd1 vssd1 vccd1 vccd1 _03234_
+ sky130_fd_sc_hd__nor2_1
XFILLER_235_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21196_ _00245_ _01212_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20147_ rbzero.texV\[-4\] _02989_ _03142_ _03176_ vssd1 vssd1 vccd1 vccd1 _01314_
+ sky130_fd_sc_hd__a22o_1
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20078_ _03130_ vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__clkinv_2
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11920_ gpout0.vpos\[0\] vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__buf_2
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11851_ rbzero.tex_b1\[30\] _03934_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__and2_1
XFILLER_79_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10802_ rbzero.tex_g0\[30\] rbzero.tex_g0\[29\] _03616_ vssd1 vssd1 vccd1 vccd1 _03625_
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ rbzero.wall_tracer.stepDistY\[9\] _07237_ _04925_ vssd1 vssd1 vccd1 vccd1
+ _07238_ sky130_fd_sc_hd__mux2_1
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11782_ _03994_ _04492_ _04496_ _03900_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__a211o_1
XFILLER_54_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13521_ _06181_ _06209_ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ _03588_ vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16240_ _08850_ vssd1 vssd1 vccd1 vccd1 _08851_ sky130_fd_sc_hd__buf_2
XFILLER_202_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ _06114_ _06119_ _06118_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__o21a_1
XFILLER_201_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10664_ rbzero.tex_g1\[31\] rbzero.tex_g1\[32\] _03552_ vssd1 vssd1 vccd1 vccd1 _03553_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12403_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__xor2_2
XFILLER_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16171_ _07229_ _08474_ _07234_ vssd1 vssd1 vccd1 vccd1 _08783_ sky130_fd_sc_hd__o21ai_1
XFILLER_167_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13383_ _05629_ _05622_ _05626_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__o21ai_1
XFILLER_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10595_ _03516_ vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15122_ _07735_ vssd1 vssd1 vccd1 vccd1 _07736_ sky130_fd_sc_hd__buf_2
X_12334_ _03798_ _04939_ _05027_ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__o21ai_4
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15053_ _07202_ _07448_ vssd1 vssd1 vccd1 vccd1 _07667_ sky130_fd_sc_hd__xnor2_2
X_19930_ _03116_ vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__clkinv_2
X_12265_ rbzero.wall_tracer.trackDistX\[2\] _04942_ rbzero.wall_tracer.trackDistX\[1\]
+ _04944_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__a22o_1
XFILLER_141_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14004_ _05638_ _06389_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__nor2_1
XFILLER_107_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11216_ _03934_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__buf_4
XFILLER_141_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19861_ _03109_ vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__clkinv_2
XFILLER_64_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12196_ net47 _04899_ _04900_ o_tex_oeb0 _04901_ vssd1 vssd1 vccd1 vccd1 _04902_
+ sky130_fd_sc_hd__a221o_1
X_18812_ _02528_ _02529_ _02530_ _02531_ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__a211o_1
XFILLER_214_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11147_ _03840_ _03865_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__or2_1
X_19792_ _04106_ _02719_ _02742_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__o21ai_1
XFILLER_228_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18743_ _02465_ _02467_ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__and2_1
XTAP_5360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15955_ _08035_ _08109_ vssd1 vssd1 vccd1 vccd1 _08569_ sky130_fd_sc_hd__or2_1
XFILLER_114_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11078_ rbzero.vga_sync.vsync _03442_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__nor2_1
XTAP_5371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14906_ _07519_ _07509_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__nor2_4
XTAP_5393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18674_ _09256_ _02403_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__nor2_1
X_15886_ _07857_ _07868_ _07856_ vssd1 vssd1 vccd1 vccd1 _08500_ sky130_fd_sc_hd__a21bo_1
XFILLER_188_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17625_ _10041_ _10160_ vssd1 vssd1 vccd1 vccd1 _10161_ sky130_fd_sc_hd__xor2_1
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14837_ _07342_ _05203_ vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__nand2_1
XFILLER_149_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17556_ _09975_ _09984_ _09983_ vssd1 vssd1 vccd1 vccd1 _10093_ sky130_fd_sc_hd__a21bo_1
XFILLER_189_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14768_ _07341_ _05091_ vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__nor2_1
XFILLER_225_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16507_ _07632_ _09115_ vssd1 vssd1 vccd1 vccd1 _09116_ sky130_fd_sc_hd__or2_1
XFILLER_220_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13719_ _05738_ _06407_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__nand2_1
XFILLER_149_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17487_ _10023_ _10024_ vssd1 vssd1 vccd1 vccd1 _10025_ sky130_fd_sc_hd__nand2_1
X_14699_ rbzero.wall_tracer.stepDistX\[4\] _07217_ _07316_ vssd1 vssd1 vccd1 vccd1
+ _07324_ sky130_fd_sc_hd__mux2_1
XFILLER_225_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19226_ _02794_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__clkbuf_4
X_16438_ _08478_ _08928_ _07826_ vssd1 vssd1 vccd1 vccd1 _09048_ sky130_fd_sc_hd__a21o_1
XFILLER_149_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19157_ rbzero.spi_registers.got_new_sky _02720_ vssd1 vssd1 vccd1 vccd1 _02752_
+ sky130_fd_sc_hd__nand2_2
X_16369_ _08978_ vssd1 vssd1 vccd1 vccd1 _08979_ sky130_fd_sc_hd__clkbuf_4
XFILLER_157_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18108_ _01853_ _01888_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__xor2_1
XFILLER_195_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19088_ _02707_ vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18039_ _01711_ _01720_ _01820_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a21oi_1
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21050_ _00099_ _01066_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20001_ _03122_ vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__clkinv_2
XFILLER_232_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20903_ net61 _00919_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20834_ _00052_ _00850_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_230_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20765_ net106 _00781_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_floor
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20696_ net99 _00712_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10380_ rbzero.tex_r1\[36\] rbzero.tex_r1\[37\] _03400_ vssd1 vssd1 vccd1 vccd1 _03402_
+ sky130_fd_sc_hd__mux2_1
XFILLER_163_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21317_ _00340_ _01333_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12050_ net47 _04748_ _04749_ net48 vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a22o_1
X_21248_ _00297_ _01264_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11001_ _03728_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__buf_4
XFILLER_46_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21179_ _00228_ _01195_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15740_ _08271_ _08314_ vssd1 vssd1 vccd1 vccd1 _08354_ sky130_fd_sc_hd__xor2_1
XFILLER_111_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _05640_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__clkbuf_4
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11903_ net13 _04612_ _04613_ net12 vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__a31o_1
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _08155_ _08282_ vssd1 vssd1 vccd1 vccd1 _08285_ sky130_fd_sc_hd__and2b_1
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _05353_ _05430_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__nor2_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _09914_ _09846_ _09946_ vssd1 vssd1 vccd1 vccd1 _09948_ sky130_fd_sc_hd__nand3_1
XFILLER_2_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ rbzero.wall_tracer.visualWallDist\[-3\] _07253_ _07276_ _07277_ _07266_ vssd1
+ vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__o221a_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ rbzero.tex_b1\[33\] rbzero.tex_b1\[32\] _04032_ vssd1 vssd1 vccd1 vccd1 _04548_
+ sky130_fd_sc_hd__mux2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ rbzero.debug_overlay.vplaneX\[-5\] rbzero.wall_tracer.rayAddendX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__nand2_1
XFILLER_92_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _09660_ _09751_ _09879_ vssd1 vssd1 vccd1 vccd1 _09880_ sky130_fd_sc_hd__a21oi_1
XFILLER_183_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14553_ _07082_ _07214_ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__or2_1
XFILLER_109_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11765_ _03956_ _04467_ _04471_ _04479_ _03985_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__o311a_1
XFILLER_199_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13504_ _06191_ _06192_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__and2_1
XFILLER_18_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10716_ rbzero.tex_g1\[6\] rbzero.tex_g1\[7\] _03574_ vssd1 vssd1 vccd1 vccd1 _03580_
+ sky130_fd_sc_hd__mux2_1
X_17272_ _08732_ _09571_ _09429_ _07618_ vssd1 vssd1 vccd1 vccd1 _09811_ sky130_fd_sc_hd__o22ai_1
X_14484_ _05527_ _07123_ _07167_ _05535_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__o211a_1
XFILLER_159_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11696_ _04410_ _04411_ _03968_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__mux2_1
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19011_ _02666_ vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16223_ _08833_ _08834_ vssd1 vssd1 vccd1 vccd1 _08835_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13435_ _06104_ _06105_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__and2_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ rbzero.tex_g1\[39\] rbzero.tex_g1\[40\] _03541_ vssd1 vssd1 vccd1 vccd1 _03544_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16154_ _08764_ _08765_ vssd1 vssd1 vccd1 vccd1 _08766_ sky130_fd_sc_hd__nand2_1
XFILLER_173_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13366_ _06053_ _06041_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__or2b_1
XFILLER_155_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10578_ _03507_ vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__clkbuf_1
X_15105_ _07670_ _07718_ vssd1 vssd1 vccd1 vccd1 _07719_ sky130_fd_sc_hd__nor2_1
X_12317_ _04961_ _04990_ _05010_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__a21oi_1
XFILLER_170_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16085_ _08589_ _08696_ vssd1 vssd1 vccd1 vccd1 _08698_ sky130_fd_sc_hd__nand2_1
XFILLER_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13297_ _05793_ _05610_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__nor2_1
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12248_ rbzero.wall_tracer.trackDistY\[2\] vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__inv_2
X_15036_ _07337_ _07649_ _07408_ vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__a21o_1
XFILLER_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19913_ _03113_ vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__clkinv_2
XFILLER_218_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19844_ _03107_ vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__clkinv_2
X_12179_ net36 net35 vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__nor2_1
XFILLER_9_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19775_ _04111_ gpout0.vpos\[6\] _04104_ _04106_ vssd1 vssd1 vccd1 vccd1 _03082_
+ sky130_fd_sc_hd__or4_1
X_16987_ _09445_ _09425_ vssd1 vssd1 vccd1 vccd1 _09528_ sky130_fd_sc_hd__or2b_1
XFILLER_228_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18726_ _02450_ _02451_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__xor2_1
X_15938_ _08550_ _08551_ vssd1 vssd1 vccd1 vccd1 _08552_ sky130_fd_sc_hd__xnor2_2
XTAP_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18657_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.wall_tracer.rayAddendY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__nand2_1
X_15869_ _08481_ _08482_ vssd1 vssd1 vccd1 vccd1 _08483_ sky130_fd_sc_hd__nor2_1
XFILLER_188_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17608_ _10143_ _10144_ vssd1 vssd1 vccd1 vccd1 _10145_ sky130_fd_sc_hd__or2b_1
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18588_ _02274_ rbzero.wall_tracer.rayAddendX\[9\] vssd1 vssd1 vccd1 vccd1 _02328_
+ sky130_fd_sc_hd__or2_1
XFILLER_224_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_150 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_150/HI o_rgb[10]
+ sky130_fd_sc_hd__conb_1
XFILLER_75_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17539_ _09571_ _08735_ _10075_ vssd1 vssd1 vccd1 vccd1 _10076_ sky130_fd_sc_hd__or3_1
XFILLER_36_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20550_ net124 _00566_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19209_ _02578_ _02784_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__or2_1
XFILLER_192_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20481_ net96 _00497_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.side sky130_fd_sc_hd__dfxtp_1
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21102_ _00151_ _01118_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout102 net104 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_236_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout113 net115 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_2
X_21033_ _00082_ _01049_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[1\] sky130_fd_sc_hd__dfxtp_1
Xfanout124 net125 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_2
Xfanout135 net139 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_2
XFILLER_160_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20817_ _00035_ _00833_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11550_ rbzero.debug_overlay.facingY\[-9\] _04240_ _04218_ rbzero.debug_overlay.facingY\[-8\]
+ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__a22o_1
XFILLER_243_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20748_ net103 _00764_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10501_ rbzero.tex_r0\[45\] rbzero.tex_r0\[44\] _03457_ vssd1 vssd1 vccd1 vccd1 _03467_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11481_ _04197_ _04198_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__or2b_1
XFILLER_17_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20679_ net76 _00695_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_183_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ _05791_ _05908_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__xor2_1
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10432_ rbzero.tex_r1\[11\] rbzero.tex_r1\[12\] _03422_ vssd1 vssd1 vccd1 vccd1 _03429_
+ sky130_fd_sc_hd__mux2_1
XFILLER_195_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13151_ _05780_ _05737_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__or2b_1
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10363_ rbzero.tex_r1\[44\] rbzero.tex_r1\[45\] _03389_ vssd1 vssd1 vccd1 vccd1 _03393_
+ sky130_fd_sc_hd__mux2_1
XFILLER_191_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12102_ _04115_ _04797_ _04809_ gpout3.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _04810_
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13082_ _05766_ _05700_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__nand2_1
XFILLER_139_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10294_ _03356_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16910_ _09449_ _09451_ _09190_ vssd1 vssd1 vccd1 vccd1 _09452_ sky130_fd_sc_hd__or3b_1
X_12033_ net5 _04738_ _04719_ _04741_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__a22o_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17890_ _01671_ _01672_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16841_ _09140_ _09154_ _09152_ vssd1 vssd1 vccd1 vccd1 _09383_ sky130_fd_sc_hd__a21o_1
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19560_ net51 rbzero.pov.ss_buffer\[0\] _02708_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__mux2_1
X_16772_ _09318_ _09319_ _09320_ vssd1 vssd1 vccd1 vccd1 _09321_ sky130_fd_sc_hd__nand3_1
XFILLER_219_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13984_ _06665_ _06666_ _06671_ vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__nand3_1
XFILLER_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18511_ _09261_ _02250_ _02251_ _02256_ vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__a31o_1
XFILLER_207_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15723_ _07789_ _07593_ _07646_ _07718_ vssd1 vssd1 vccd1 vccd1 _08337_ sky130_fd_sc_hd__or4_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12935_ _05582_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__clkbuf_4
X_19491_ _02913_ vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18442_ _02191_ rbzero.wall_tracer.rayAddendX\[-1\] vssd1 vssd1 vccd1 vccd1 _02192_
+ sky130_fd_sc_hd__nand2_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _08248_ _08266_ vssd1 vssd1 vccd1 vccd1 _08268_ sky130_fd_sc_hd__or2b_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12866_ _05497_ _05456_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__nor2_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _03819_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__clkbuf_4
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18373_ _01823_ _02130_ _01996_ rbzero.wall_tracer.trackDistY\[9\] vssd1 vssd1 vccd1
+ vccd1 _00586_ sky130_fd_sc_hd__o2bb2a_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ rbzero.tex_b1\[58\] _03934_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__and2_1
X_15585_ _07481_ _07482_ _07483_ _07645_ vssd1 vssd1 vccd1 vccd1 _08199_ sky130_fd_sc_hd__a211o_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12797_ _05484_ _05485_ _05453_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__mux2_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17324_ _09859_ _09860_ _09862_ vssd1 vssd1 vccd1 vccd1 _09863_ sky130_fd_sc_hd__and3_1
XFILLER_42_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14536_ _07133_ _07052_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__or2_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11748_ _03994_ _04458_ _04462_ _03900_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__a211o_1
XFILLER_239_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17255_ _09792_ _09793_ vssd1 vssd1 vccd1 vccd1 _09794_ sky130_fd_sc_hd__or2b_1
X_14467_ _07105_ _07125_ _07152_ _07107_ vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__a211o_1
XFILLER_128_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11679_ _04392_ _04393_ _04394_ _03958_ _03994_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__o221a_1
X_16206_ _08814_ _08816_ vssd1 vssd1 vccd1 vccd1 _08818_ sky130_fd_sc_hd__nand2_1
XFILLER_128_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13418_ _05793_ _05635_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__nor2_1
XFILLER_31_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17186_ _09719_ _09725_ vssd1 vssd1 vccd1 vccd1 _09726_ sky130_fd_sc_hd__xnor2_1
XFILLER_122_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14398_ _07029_ _07060_ vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__or2_1
XFILLER_196_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16137_ _07469_ _08274_ _08067_ _07790_ vssd1 vssd1 vccd1 vccd1 _08749_ sky130_fd_sc_hd__or4_1
XFILLER_155_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13349_ _05997_ _06014_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__xor2_1
XFILLER_127_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16068_ _08534_ _08543_ _08541_ vssd1 vssd1 vccd1 vccd1 _08681_ sky130_fd_sc_hd__o21a_1
XFILLER_170_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15019_ _03794_ rbzero.wall_tracer.stepDistY\[-12\] _07632_ vssd1 vssd1 vccd1 vccd1
+ _07633_ sky130_fd_sc_hd__o21ai_4
XFILLER_237_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19827_ _03106_ vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__clkinv_2
XFILLER_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19758_ rbzero.pov.ready_buffer\[8\] _03055_ _03058_ rbzero.debug_overlay.vplaneY\[-1\]
+ _02832_ vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__o221a_1
XFILLER_186_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18709_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.debug_overlay.vplaneY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__nor2_1
XFILLER_204_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19689_ rbzero.pov.ready_buffer\[56\] _02963_ _03044_ _03045_ _03012_ vssd1 vssd1
+ vccd1 vccd1 _03046_ sky130_fd_sc_hd__o221a_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20602_ net82 _00618_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_240_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20533_ net123 _00549_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20464_ net118 _00480_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.side sky130_fd_sc_hd__dfxtp_2
XFILLER_14_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20395_ net137 _00426_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21016_ net57 _01032_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_5937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10981_ rbzero.tex_b0\[9\] rbzero.tex_b0\[8\] _03715_ vssd1 vssd1 vccd1 vccd1 _03719_
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12720_ _05373_ _05361_ _05363_ _05375_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__or4b_1
XFILLER_16_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12651_ _05211_ _05213_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__nand2_2
XFILLER_231_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ rbzero.tex_g0\[3\] _03939_ _03941_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__and3_1
X_15370_ _04935_ rbzero.wall_tracer.stepDistX\[-11\] vssd1 vssd1 vccd1 vccd1 _07984_
+ sky130_fd_sc_hd__nand2_1
X_12582_ _05265_ _05270_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__nand2b_1
XFILLER_230_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14321_ _07008_ _07009_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__or2_1
XFILLER_157_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11533_ rbzero.debug_overlay.facingX\[-3\] _04209_ _04219_ _04250_ vssd1 vssd1 vccd1
+ vccd1 _04251_ sky130_fd_sc_hd__a211o_1
XFILLER_180_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17040_ _09172_ _09434_ _09436_ _09437_ vssd1 vssd1 vccd1 vccd1 _09581_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14252_ _06921_ _06929_ vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__or2_1
X_11464_ _03924_ _04177_ _04181_ _03950_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__a211o_1
XFILLER_137_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13203_ _05890_ _05891_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__xnor2_1
X_10415_ rbzero.tex_r1\[19\] rbzero.tex_r1\[20\] _03411_ vssd1 vssd1 vccd1 vccd1 _03420_
+ sky130_fd_sc_hd__mux2_1
XFILLER_165_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14183_ _06870_ _06871_ vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__nor2_1
XFILLER_139_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11395_ _04104_ _04113_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__nand2_1
XFILLER_178_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13134_ _05699_ _05700_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__nand2_1
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10346_ _03383_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__clkbuf_1
X_18991_ rbzero.pov.spi_buffer\[43\] rbzero.pov.ready_buffer\[43\] _02651_ vssd1 vssd1
+ vccd1 vccd1 _02656_ sky130_fd_sc_hd__mux2_1
XFILLER_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17942_ _01613_ _01615_ _01614_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__a21boi_1
X_13065_ _05744_ _05753_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10277_ _03347_ vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12016_ _04717_ o_rgb[7] _04724_ net7 vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__a211o_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17873_ _01654_ _01655_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__xor2_1
XFILLER_79_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16824_ _07332_ _09365_ _09366_ _09275_ vssd1 vssd1 vccd1 vccd1 _09367_ sky130_fd_sc_hd__o31a_1
X_19612_ rbzero.debug_overlay.playerX\[1\] _02982_ _02962_ vssd1 vssd1 vccd1 vccd1
+ _02986_ sky130_fd_sc_hd__o21ai_1
XFILLER_120_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19543_ _02940_ vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16755_ _09295_ _09296_ _09297_ vssd1 vssd1 vccd1 vccd1 _09306_ sky130_fd_sc_hd__o21bai_1
XFILLER_150_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13967_ _06646_ _06647_ _06655_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15706_ _08315_ _08317_ vssd1 vssd1 vccd1 vccd1 _08320_ sky130_fd_sc_hd__nor2_1
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12918_ _05537_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__buf_2
XFILLER_62_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19474_ _02904_ vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__clkbuf_1
XFILLER_222_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16686_ rbzero.traced_texa\[-10\] _09262_ _09263_ rbzero.wall_tracer.visualWallDist\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__a22o_1
XFILLER_59_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13898_ _06510_ _06586_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__nand2_1
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18425_ _02174_ _02176_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__xnor2_1
XFILLER_206_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15637_ _08227_ _08226_ vssd1 vssd1 vccd1 vccd1 _08251_ sky130_fd_sc_hd__xor2_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12849_ _05440_ _05470_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__nor2_2
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18356_ _02113_ _02114_ _02115_ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__a21oi_1
XFILLER_194_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15568_ _07377_ _07398_ _07507_ _07592_ vssd1 vssd1 vccd1 vccd1 _08182_ sky130_fd_sc_hd__or4_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17307_ _09826_ _09845_ vssd1 vssd1 vccd1 vccd1 _09846_ sky130_fd_sc_hd__nand2_1
XFILLER_187_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14519_ _07197_ vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18287_ _09345_ _02055_ _02056_ _09352_ _01995_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__o311a_1
X_15499_ _08104_ _08101_ vssd1 vssd1 vccd1 vccd1 _08113_ sky130_fd_sc_hd__and2b_1
XFILLER_174_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17238_ _09662_ _09695_ vssd1 vssd1 vccd1 vccd1 _09777_ sky130_fd_sc_hd__nand2_1
XFILLER_163_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17169_ _08760_ _08628_ vssd1 vssd1 vccd1 vccd1 _09709_ sky130_fd_sc_hd__nor2_1
XFILLER_31_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20180_ _03093_ _03203_ _03204_ _03064_ rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1
+ _01319_ sky130_fd_sc_hd__a32o_1
XFILLER_143_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20516_ net132 _00532_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20447_ net95 _00013_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10200_ rbzero.tex_b1\[57\] rbzero.tex_b1\[58\] _03300_ vssd1 vssd1 vccd1 vccd1 _03307_
+ sky130_fd_sc_hd__mux2_1
XFILLER_106_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11180_ _03898_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__buf_4
XFILLER_101_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20378_ net116 _00409_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_7136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14870_ _07481_ _07482_ _07483_ vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__a21o_1
XFILLER_134_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13821_ _05641_ _06320_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__nand2_2
XFILLER_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16540_ _09141_ _09148_ vssd1 vssd1 vccd1 vccd1 _09149_ sky130_fd_sc_hd__xnor2_1
XFILLER_216_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13752_ _05740_ _06312_ _06440_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__o21ai_1
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10964_ rbzero.tex_b0\[17\] rbzero.tex_b0\[16\] _03704_ vssd1 vssd1 vccd1 vccd1 _03710_
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12703_ _05322_ _05383_ _05388_ _05390_ _05391_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__a41o_1
XFILLER_56_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16471_ _09077_ _09078_ _09080_ vssd1 vssd1 vccd1 vccd1 _09081_ sky130_fd_sc_hd__nand3_1
X_13683_ _06351_ _06360_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10895_ rbzero.tex_b0\[50\] rbzero.tex_b0\[49\] _03671_ vssd1 vssd1 vccd1 vccd1 _03674_
+ sky130_fd_sc_hd__mux2_1
X_18210_ _05121_ _01988_ _01989_ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__or3b_2
XFILLER_223_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15422_ _08002_ _08032_ vssd1 vssd1 vccd1 vccd1 _08036_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12634_ _05311_ _05316_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__xnor2_2
X_19190_ rbzero.spi_registers.got_new_vshift _02721_ vssd1 vssd1 vccd1 vccd1 _02773_
+ sky130_fd_sc_hd__and2_1
XFILLER_93_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18141_ _01916_ _01921_ rbzero.wall_tracer.trackDistX\[10\] _09276_ vssd1 vssd1 vccd1
+ vccd1 _00563_ sky130_fd_sc_hd__o2bb2a_1
X_15353_ _07378_ _07399_ _07423_ _07485_ vssd1 vssd1 vccd1 vccd1 _07967_ sky130_fd_sc_hd__nor4_1
XFILLER_145_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12565_ rbzero.wall_tracer.visualWallDist\[-11\] rbzero.wall_tracer.rayAddendY\[-3\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__mux2_1
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14304_ _06455_ _06974_ vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__xor2_1
X_18072_ _01835_ _01852_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__xnor2_1
X_11516_ _04232_ _04233_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__and2_1
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15284_ _07896_ _07897_ vssd1 vssd1 vccd1 vccd1 _07898_ sky130_fd_sc_hd__and2b_1
XFILLER_184_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12496_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[11\] vssd1
+ vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__nor2_2
XFILLER_172_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17023_ _09443_ _09528_ _09562_ vssd1 vssd1 vccd1 vccd1 _09564_ sky130_fd_sc_hd__and3_1
X_14235_ _06913_ _06918_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11447_ rbzero.tex_r1\[27\] rbzero.tex_r1\[26\] _03904_ vssd1 vssd1 vccd1 vccd1 _04165_
+ sky130_fd_sc_hd__mux2_1
XFILLER_236_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14166_ _06851_ _06854_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__and2_1
X_11378_ rbzero.row_render.size\[10\] rbzero.row_render.size\[9\] _04047_ _04096_
+ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__or4_2
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13117_ _05804_ _05805_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__xnor2_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _03374_ vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__clkbuf_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _06783_ _06784_ _06785_ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__a21oi_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18974_ rbzero.pov.spi_buffer\[35\] rbzero.pov.ready_buffer\[35\] _02640_ vssd1 vssd1
+ vccd1 vccd1 _02647_ sky130_fd_sc_hd__mux2_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ _01705_ _01707_ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__xnor2_1
X_13048_ _05698_ _05735_ _05736_ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__o21ai_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17856_ _09968_ _09603_ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__nor2_1
XFILLER_120_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16807_ _09351_ _08959_ vssd1 vssd1 vccd1 vccd1 _09352_ sky130_fd_sc_hd__nand2_1
XFILLER_113_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17787_ _07631_ _07827_ _01570_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__or3_1
X_14999_ _07605_ _07611_ vssd1 vssd1 vccd1 vccd1 _07613_ sky130_fd_sc_hd__nor2_1
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16738_ _09279_ _09289_ _09290_ _09283_ vssd1 vssd1 vccd1 vccd1 _09291_ sky130_fd_sc_hd__a31o_1
X_19526_ _02931_ vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_223_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19457_ _02895_ vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__clkbuf_1
X_16669_ rbzero.row_render.size\[6\] _09255_ _07196_ _09259_ vssd1 vssd1 vccd1 vccd1
+ _00504_ sky130_fd_sc_hd__a22o_1
XFILLER_35_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18408_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__and2_1
X_19388_ _02861_ vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__clkinv_2
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18339_ rbzero.wall_tracer.trackDistY\[5\] rbzero.wall_tracer.stepDistY\[5\] vssd1
+ vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__nor2_1
XFILLER_202_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21350_ _00373_ _01366_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20301_ _03258_ vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__clkinv_2
X_21281_ _00330_ _01297_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20232_ _03245_ _03246_ _03247_ _03240_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__a22o_1
XFILLER_196_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20163_ _03183_ _03187_ _03188_ _03189_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__o211a_1
XFILLER_157_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20094_ gpout5.clk_div\[1\] gpout5.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__or2_1
XFILLER_69_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20996_ net55 _01012_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10680_ rbzero.tex_g1\[23\] rbzero.tex_g1\[24\] _03552_ vssd1 vssd1 vccd1 vccd1 _03561_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12350_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] _05038_
+ _05041_ _05042_ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__a221o_1
XFILLER_217_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11301_ _04018_ _04019_ _03932_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__mux2_1
XFILLER_181_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12281_ _04964_ _04974_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__nor2_1
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14020_ _06706_ _06708_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__nor2_1
XFILLER_135_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11232_ _03924_ _03931_ _03947_ _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__a211o_1
XFILLER_135_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11163_ rbzero.traced_texVinit\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _03882_
+ sky130_fd_sc_hd__xnor2_1
XTAP_6210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15971_ _07334_ _05114_ _08584_ vssd1 vssd1 vccd1 vccd1 _08585_ sky130_fd_sc_hd__o21ai_4
X_11094_ _03792_ _03729_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__nor2_1
XFILLER_49_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17710_ _10047_ _10138_ _10136_ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__a21oi_1
XTAP_6287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14922_ rbzero.wall_tracer.visualWallDist\[-3\] _07535_ _07349_ vssd1 vssd1 vccd1
+ vccd1 _07536_ sky130_fd_sc_hd__mux2_1
XFILLER_236_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18690_ _04260_ rbzero.wall_tracer.rayAddendY\[-2\] _02410_ vssd1 vssd1 vccd1 vccd1
+ _02418_ sky130_fd_sc_hd__a21o_1
XFILLER_236_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17641_ _01424_ _01425_ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__and2_1
XTAP_5597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14853_ _07460_ _07461_ _07465_ _07466_ vssd1 vssd1 vccd1 vccd1 _07467_ sky130_fd_sc_hd__a22o_2
XFILLER_76_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13804_ _06460_ _06466_ _06492_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__o21a_1
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17572_ _10092_ _10108_ vssd1 vssd1 vccd1 vccd1 _10109_ sky130_fd_sc_hd__xnor2_1
X_14784_ _07356_ _07392_ _07393_ _07397_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__o31ai_4
XFILLER_205_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11996_ net48 _04664_ net15 vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__and3_1
XFILLER_204_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19311_ _02845_ vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__clkbuf_1
X_16523_ _09130_ _09131_ vssd1 vssd1 vccd1 vccd1 _09132_ sky130_fd_sc_hd__and2b_1
XFILLER_204_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13735_ _05861_ _06423_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__or2_1
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10947_ rbzero.tex_b0\[25\] rbzero.tex_b0\[24\] _03693_ vssd1 vssd1 vccd1 vccd1 _03701_
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19242_ _02803_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__buf_2
X_16454_ _09059_ _09060_ _09062_ vssd1 vssd1 vccd1 vccd1 _09064_ sky130_fd_sc_hd__a21o_1
XFILLER_220_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13666_ _06353_ _06354_ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__and2b_1
XFILLER_147_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10878_ rbzero.tex_b0\[58\] rbzero.tex_b0\[57\] _03660_ vssd1 vssd1 vccd1 vccd1 _03665_
+ sky130_fd_sc_hd__mux2_1
XFILLER_188_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15405_ _07945_ _08006_ _08018_ vssd1 vssd1 vccd1 vccd1 _08019_ sky130_fd_sc_hd__a21o_1
XFILLER_160_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _05277_ _05289_ _05304_ _05305_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__o31a_1
X_19173_ _02762_ vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__clkbuf_1
X_16385_ _08866_ _08868_ _08865_ vssd1 vssd1 vccd1 vccd1 _08995_ sky130_fd_sc_hd__a21bo_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ _06263_ _06284_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__nor2_1
XFILLER_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18124_ _01901_ _01903_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__nand2_1
XFILLER_160_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15336_ _07947_ _07948_ _07949_ vssd1 vssd1 vccd1 vccd1 _07950_ sky130_fd_sc_hd__a21oi_1
X_12548_ _05219_ _05236_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__or2_1
XFILLER_247_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18055_ _01746_ _01747_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__or2_1
X_15267_ _07485_ _07591_ _07790_ _07880_ vssd1 vssd1 vccd1 vccd1 _07881_ sky130_fd_sc_hd__or4_1
XANTENNA_2 _01823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _05155_ _05158_ _05164_ _05167_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__and4bb_1
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17006_ _09430_ _09432_ _09427_ vssd1 vssd1 vccd1 vccd1 _09547_ sky130_fd_sc_hd__a21bo_1
X_14218_ _06899_ _06900_ vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__or2_1
XFILLER_119_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15198_ _07784_ _07811_ vssd1 vssd1 vccd1 vccd1 _07812_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14149_ _06809_ _06835_ _06837_ vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__and3_1
XFILLER_119_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18957_ rbzero.pov.spi_buffer\[27\] rbzero.pov.ready_buffer\[27\] _02629_ vssd1 vssd1
+ vccd1 vccd1 _02638_ sky130_fd_sc_hd__mux2_1
XFILLER_112_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17908_ _01562_ _01527_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__or2b_1
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18888_ _02599_ vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17839_ _10121_ _01621_ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__xor2_1
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20850_ _00068_ _00866_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19509_ rbzero.pov.spi_buffer\[50\] rbzero.pov.spi_buffer\[51\] _02921_ vssd1 vssd1
+ vccd1 vccd1 _02923_ sky130_fd_sc_hd__mux2_1
XFILLER_212_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20781_ net87 _00797_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21402_ net110 _01418_ vssd1 vssd1 vccd1 vccd1 gpout2.clk_div\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21333_ _00356_ _01349_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21264_ _00313_ _01280_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20215_ rbzero.texV\[7\] _03137_ _03142_ _03233_ vssd1 vssd1 vccd1 vccd1 _01325_
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21195_ _00244_ _01211_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20146_ _03173_ _03175_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__xnor2_1
XFILLER_132_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20077_ _03130_ vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__clkinv_2
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ rbzero.tex_b1\[29\] rbzero.tex_b1\[28\] _03934_ vssd1 vssd1 vccd1 vccd1 _04564_
+ sky130_fd_sc_hd__mux2_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10801_ _03624_ vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__clkbuf_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11781_ _04323_ _04493_ _04494_ _04495_ _03921_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__o221a_1
XFILLER_72_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20979_ net65 _00995_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13520_ _06193_ _06208_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__xnor2_1
XFILLER_242_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10732_ rbzero.tex_g0\[63\] rbzero.tex_g0\[62\] _03512_ vssd1 vssd1 vccd1 vccd1 _03588_
+ sky130_fd_sc_hd__mux2_1
XFILLER_246_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13451_ _06136_ _06138_ _06139_ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__or3_1
XFILLER_90_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10663_ _03388_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__clkbuf_4
XFILLER_220_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12402_ _05094_ _05039_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__xnor2_2
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16170_ _07229_ _07234_ _08474_ vssd1 vssd1 vccd1 vccd1 _08782_ sky130_fd_sc_hd__or3_1
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13382_ _05629_ _05715_ _05626_ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__or3_1
XFILLER_51_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10594_ rbzero.tex_r0\[1\] rbzero.tex_r0\[0\] _03512_ vssd1 vssd1 vccd1 vccd1 _03516_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15121_ _04935_ _07729_ _07733_ _07734_ vssd1 vssd1 vccd1 vccd1 _07735_ sky130_fd_sc_hd__o31a_2
XFILLER_127_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12333_ _04940_ _05025_ _05026_ vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__o21a_2
XFILLER_103_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15052_ _07654_ _07665_ vssd1 vssd1 vccd1 vccd1 _07666_ sky130_fd_sc_hd__xor2_1
XFILLER_114_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12264_ _04952_ _04955_ _04956_ _04957_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__a211o_1
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14003_ _05740_ _06343_ _06305_ _06028_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__a2bb2o_1
X_11215_ _03902_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__clkbuf_4
X_12195_ net48 net34 _04874_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__and3_1
X_19860_ _03109_ vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__clkinv_2
X_18811_ rbzero.wall_tracer.rayAddendY\[6\] rbzero.wall_tracer.rayAddendY\[5\] rbzero.wall_tracer.rayAddendY\[4\]
+ rbzero.wall_tracer.rayAddendY\[3\] _02509_ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__o41a_1
XFILLER_110_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11146_ _03836_ _03839_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__and2_1
XTAP_6051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19791_ _04106_ _03808_ _02718_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__and3_1
XTAP_6062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11077_ _03796_ _03800_ _03730_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__a21oi_1
X_15954_ _08171_ _08457_ _08169_ vssd1 vssd1 vccd1 vccd1 _08568_ sky130_fd_sc_hd__a21boi_2
X_18742_ _02448_ _02449_ _02451_ _02466_ _02436_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__a32o_1
XFILLER_231_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14905_ _04937_ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__buf_4
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18673_ _02400_ _02402_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__xnor2_1
X_15885_ _08496_ _08497_ _08471_ vssd1 vssd1 vccd1 vccd1 _08499_ sky130_fd_sc_hd__a21o_1
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17624_ _10158_ _10159_ vssd1 vssd1 vccd1 vccd1 _10160_ sky130_fd_sc_hd__nor2_1
X_14836_ _07445_ _07449_ _07337_ vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__a21oi_2
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _09960_ _09970_ _10091_ vssd1 vssd1 vccd1 vccd1 _10092_ sky130_fd_sc_hd__a21o_1
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14767_ _07213_ _07184_ _07336_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__a21o_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11979_ _04665_ _04118_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__nor2_1
XFILLER_189_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16506_ _09114_ vssd1 vssd1 vccd1 vccd1 _09115_ sky130_fd_sc_hd__clkbuf_4
XFILLER_204_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13718_ _06406_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__clkbuf_2
XFILLER_147_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17486_ _09758_ _09884_ _09883_ vssd1 vssd1 vccd1 vccd1 _10024_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14698_ _07323_ vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16437_ _07824_ _08793_ _07468_ vssd1 vssd1 vccd1 vccd1 _09047_ sky130_fd_sc_hd__a21o_1
X_19225_ _02784_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__or3b_1
X_13649_ _06337_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__inv_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19156_ rbzero.floor_leak\[5\] _02744_ _02751_ _02738_ vssd1 vssd1 vccd1 vccd1 _00748_
+ sky130_fd_sc_hd__o211a_1
X_16368_ _05301_ _08629_ _04939_ vssd1 vssd1 vccd1 vccd1 _08978_ sky130_fd_sc_hd__or3_4
XFILLER_121_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18107_ _01854_ _01887_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__xnor2_1
X_15319_ _07764_ _07770_ vssd1 vssd1 vccd1 vccd1 _07933_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19087_ rbzero.spi_registers.spi_cmd\[2\] rbzero.spi_registers.spi_cmd\[3\] _02703_
+ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__mux2_1
X_16299_ _08786_ _08790_ _08909_ vssd1 vssd1 vccd1 vccd1 _08910_ sky130_fd_sc_hd__a21o_1
XFILLER_195_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18038_ _01818_ _01819_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__or2_1
XFILLER_172_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20000_ _03122_ vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__clkinv_2
XFILLER_113_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19989_ _03121_ vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__clkinv_2
XFILLER_154_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20902_ net60 _00918_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20833_ _00051_ _00849_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20764_ net105 _00780_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20695_ net99 _00711_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_196_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21316_ _00339_ _01332_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21247_ _00296_ _01263_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11000_ o_vsync _03292_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__nand2_1
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21178_ _00227_ _01194_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20129_ _03158_ _03159_ _03160_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a21o_1
XFILLER_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _05613_ _05545_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _04611_ _04447_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__nand2_1
X_15670_ _08247_ _08267_ vssd1 vssd1 vccd1 vccd1 _08284_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _05418_ _05362_ _05463_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__mux2_1
XFILLER_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14621_ _04947_ _07246_ _07249_ vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__o21ai_1
XFILLER_27_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11833_ _04545_ _04546_ _03928_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__mux2_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _09748_ _09750_ vssd1 vssd1 vccd1 vccd1 _09879_ sky130_fd_sc_hd__nor2_1
XFILLER_187_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _06990_ _06986_ _06989_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__nand3_1
XFILLER_159_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _03924_ _04474_ _04478_ _03899_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__a211o_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13503_ _06182_ _06190_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__or2_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _07618_ _08732_ _09571_ _09429_ vssd1 vssd1 vccd1 vccd1 _09810_ sky130_fd_sc_hd__or4_1
XFILLER_41_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _03579_ vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__clkbuf_1
X_14483_ _07126_ _07128_ _07107_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__a21o_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11695_ rbzero.tex_g1\[61\] rbzero.tex_g1\[60\] _04378_ vssd1 vssd1 vccd1 vccd1 _04411_
+ sky130_fd_sc_hd__mux2_1
X_19010_ rbzero.pov.spi_buffer\[52\] rbzero.pov.ready_buffer\[52\] _02662_ vssd1 vssd1
+ vccd1 vccd1 _02666_ sky130_fd_sc_hd__mux2_1
XFILLER_109_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16222_ _08704_ _08705_ _08702_ vssd1 vssd1 vccd1 vccd1 _08834_ sky130_fd_sc_hd__o21ba_1
X_13434_ _05793_ _05671_ _05740_ _06122_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__or4_1
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10646_ _03543_ vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16153_ _08748_ _08624_ _08763_ vssd1 vssd1 vccd1 vccd1 _08765_ sky130_fd_sc_hd__nand3_1
XFILLER_31_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13365_ _06041_ _06053_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__xor2_1
XFILLER_10_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10577_ rbzero.tex_r0\[9\] rbzero.tex_r0\[8\] _03501_ vssd1 vssd1 vccd1 vccd1 _03507_
+ sky130_fd_sc_hd__mux2_1
X_15104_ _04927_ _07652_ vssd1 vssd1 vccd1 vccd1 _07718_ sky130_fd_sc_hd__nand2_2
X_12316_ _04997_ _04998_ _05000_ _05009_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__or4_1
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16084_ _08589_ _08696_ vssd1 vssd1 vccd1 vccd1 _08697_ sky130_fd_sc_hd__or2_1
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13296_ _05699_ _05567_ _05748_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__and3_1
XFILLER_138_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15035_ _05106_ _05273_ _07342_ vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__mux2_1
XFILLER_142_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19912_ _03113_ vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__clkinv_2
X_12247_ rbzero.wall_tracer.trackDistY\[3\] vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__inv_2
XFILLER_244_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19843_ _03107_ vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__clkinv_2
XFILLER_218_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12178_ _04078_ _03781_ _03784_ _03291_ _04883_ _04873_ vssd1 vssd1 vccd1 vccd1 _04884_
+ sky130_fd_sc_hd__mux4_1
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11129_ rbzero.texV\[4\] _03847_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__xor2_1
X_19774_ o_hsync _03079_ _03081_ vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__a21boi_1
XFILLER_84_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16986_ _09401_ _09402_ _09418_ _09416_ vssd1 vssd1 vccd1 vccd1 _09527_ sky130_fd_sc_hd__a31o_1
XFILLER_77_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18725_ _02422_ _02435_ _02436_ _02440_ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__o31ai_1
X_15937_ _07628_ _07921_ vssd1 vssd1 vccd1 vccd1 _08551_ sky130_fd_sc_hd__nor2_1
XTAP_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15868_ _08479_ _08480_ _08472_ vssd1 vssd1 vccd1 vccd1 _08482_ sky130_fd_sc_hd__a21oi_1
X_18656_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.wall_tracer.rayAddendY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__and2_1
XFILLER_97_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17607_ _10036_ _10037_ _10142_ vssd1 vssd1 vccd1 vccd1 _10144_ sky130_fd_sc_hd__nand3_1
XFILLER_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14819_ _07431_ _07432_ _07374_ vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__mux2_1
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15799_ _08351_ _08412_ vssd1 vssd1 vccd1 vccd1 _08413_ sky130_fd_sc_hd__nand2_1
X_18587_ _02275_ rbzero.wall_tracer.rayAddendX\[9\] vssd1 vssd1 vccd1 vccd1 _02327_
+ sky130_fd_sc_hd__nand2_1
XFILLER_18_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_151 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_151/HI o_rgb[11]
+ sky130_fd_sc_hd__conb_1
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17538_ _10073_ _10074_ vssd1 vssd1 vccd1 vccd1 _10075_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17469_ _09825_ _09873_ _10006_ vssd1 vssd1 vccd1 vccd1 _10007_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19208_ rbzero.spi_registers.spi_cmd\[3\] rbzero.spi_registers.spi_cmd\[2\] _03442_
+ rbzero.spi_registers.spi_done vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__or4b_1
X_20480_ net94 _00496_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_203_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19139_ rbzero.spi_registers.got_new_vinf _02724_ rbzero.row_render.vinf vssd1 vssd1
+ vccd1 vccd1 _02741_ sky130_fd_sc_hd__a21o_1
XFILLER_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21101_ _00150_ _01117_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_218_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21032_ _00081_ _01048_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[0\] sky130_fd_sc_hd__dfxtp_1
Xfanout103 net104 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_2
XFILLER_232_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout114 net115 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__buf_2
XFILLER_236_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout125 net126 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_113_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout136 net139 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_2
XFILLER_87_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20816_ _00034_ _00832_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20747_ net103 _00763_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_243_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10500_ _03466_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__clkbuf_1
XFILLER_149_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11480_ gpout0.hpos\[3\] _03804_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20678_ net67 _00694_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10431_ _03428_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13150_ _05784_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__nor2b_1
XFILLER_170_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10362_ _03392_ vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12101_ net26 net25 vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__nor2_1
XFILLER_30_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13081_ _05525_ _05701_ _05731_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__and3_1
X_10293_ rbzero.tex_b1\[13\] rbzero.tex_b1\[14\] _03355_ vssd1 vssd1 vccd1 vccd1 _03356_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12032_ _04739_ _04740_ _04718_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__mux2_1
XFILLER_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ _09371_ _09381_ vssd1 vssd1 vccd1 vccd1 _09382_ sky130_fd_sc_hd__xor2_1
XFILLER_215_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16771_ _09311_ _09313_ _09312_ vssd1 vssd1 vccd1 vccd1 _09320_ sky130_fd_sc_hd__o21bai_1
XFILLER_111_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13983_ _06665_ _06666_ _06671_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__a21o_1
XFILLER_150_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15722_ _07593_ _07646_ _08335_ _07789_ vssd1 vssd1 vccd1 vccd1 _08336_ sky130_fd_sc_hd__o22a_1
X_18510_ rbzero.wall_tracer.rayAddendX\[3\] _02197_ _02255_ _02157_ vssd1 vssd1 vccd1
+ vccd1 _02256_ sky130_fd_sc_hd__a22o_1
X_12934_ _05621_ _05622_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__or2_1
XFILLER_111_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19490_ rbzero.pov.spi_buffer\[41\] rbzero.pov.spi_buffer\[42\] _02910_ vssd1 vssd1
+ vccd1 vccd1 _02913_ sky130_fd_sc_hd__mux2_1
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15653_ _08248_ _08266_ vssd1 vssd1 vccd1 vccd1 _08267_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18441_ rbzero.debug_overlay.vplaneX\[-1\] vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__buf_2
XFILLER_185_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12865_ _05318_ _05321_ _05430_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__mux2_1
XFILLER_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _04963_ _07246_ _07249_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _02128_ _02129_ _02039_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__o21a_1
XFILLER_178_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ rbzero.tex_b1\[57\] rbzero.tex_b1\[56\] _04032_ vssd1 vssd1 vccd1 vccd1 _04530_
+ sky130_fd_sc_hd__mux2_1
X_15584_ _08139_ _08197_ vssd1 vssd1 vccd1 vccd1 _08198_ sky130_fd_sc_hd__xor2_2
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _05325_ _05327_ _05448_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__mux2_1
XFILLER_57_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _09730_ _09735_ _09861_ vssd1 vssd1 vccd1 vccd1 _09862_ sky130_fd_sc_hd__a21o_1
XFILLER_226_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14535_ _07209_ vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11747_ _04459_ _04460_ _04461_ _03958_ _03924_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__o221a_1
XFILLER_187_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17254_ _08596_ _08599_ _08851_ _08979_ vssd1 vssd1 vccd1 vccd1 _09793_ sky130_fd_sc_hd__or4_1
XFILLER_169_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14466_ _07105_ _07131_ vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__nor2_1
XFILLER_105_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11678_ rbzero.tex_g1\[1\] rbzero.tex_g1\[0\] _03962_ vssd1 vssd1 vccd1 vccd1 _04394_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16205_ _08814_ _08816_ vssd1 vssd1 vccd1 vccd1 _08817_ sky130_fd_sc_hd__or2_1
XFILLER_122_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13417_ _06077_ _06078_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17185_ _09723_ _09724_ vssd1 vssd1 vccd1 vccd1 _09725_ sky130_fd_sc_hd__xor2_1
XFILLER_174_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10629_ _03534_ vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__clkbuf_1
X_14397_ _05569_ _07085_ vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__nor2_1
XFILLER_183_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16136_ _08616_ _08622_ vssd1 vssd1 vccd1 vccd1 _08748_ sky130_fd_sc_hd__nand2_1
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13348_ _06029_ _06036_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__xor2_1
XFILLER_128_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16067_ _08667_ _08679_ vssd1 vssd1 vccd1 vccd1 _08680_ sky130_fd_sc_hd__xnor2_1
X_13279_ _05956_ _05961_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__o21ba_1
XFILLER_142_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15018_ _07599_ _07601_ _07352_ vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__a21oi_4
XFILLER_29_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19826_ _02862_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__buf_4
XFILLER_233_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19757_ rbzero.pov.ready_buffer\[7\] _03067_ _03068_ _04260_ _03015_ vssd1 vssd1
+ vccd1 vccd1 _01030_ sky130_fd_sc_hd__a221o_1
XFILLER_244_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16969_ _09363_ _09366_ _09509_ _09510_ vssd1 vssd1 vccd1 vccd1 _09511_ sky130_fd_sc_hd__o211a_1
XFILLER_133_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18708_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.debug_overlay.vplaneY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__and2_1
XFILLER_42_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19688_ rbzero.debug_overlay.playerY\[3\] _03039_ _02835_ vssd1 vssd1 vccd1 vccd1
+ _03045_ sky130_fd_sc_hd__a21o_1
XFILLER_224_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18639_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.wall_tracer.rayAddendY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__nor2_1
XFILLER_92_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20601_ net81 _00617_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_220_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20532_ net121 _00548_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20463_ net96 _00479_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.wall\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20394_ net138 _00425_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21015_ net57 _01031_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_5938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10980_ _03718_ vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12650_ _05220_ _05221_ _05223_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__o21ai_4
XFILLER_130_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11601_ _03899_ _04309_ _04317_ _03954_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__o211a_1
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12581_ _05220_ _05267_ _05268_ _05269_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_24_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14320_ _06962_ _06964_ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__nor2_1
XFILLER_196_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11532_ rbzero.debug_overlay.facingX\[10\] _04236_ _04239_ _04249_ vssd1 vssd1 vccd1
+ vccd1 _04250_ sky130_fd_sc_hd__a211o_1
XFILLER_19_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ _06933_ _06939_ vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__or2_1
XFILLER_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11463_ _03957_ _04178_ _04179_ _04180_ _03946_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__o221a_1
X_13202_ _05803_ _05806_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__xor2_1
XFILLER_171_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10414_ _03419_ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__clkbuf_1
X_14182_ _06869_ _06868_ vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__and2b_1
XFILLER_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11394_ _04112_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__clkbuf_2
XFILLER_109_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13133_ _05705_ _05819_ _05820_ _05821_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__o22a_1
XFILLER_125_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10345_ rbzero.tex_r1\[52\] rbzero.tex_r1\[53\] _03377_ vssd1 vssd1 vccd1 vccd1 _03383_
+ sky130_fd_sc_hd__mux2_1
X_18990_ _02655_ vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17941_ _01722_ _01723_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__and2b_1
X_13064_ _05751_ _05752_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10276_ rbzero.tex_b1\[21\] rbzero.tex_b1\[22\] _03344_ vssd1 vssd1 vccd1 vccd1 _03347_
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12015_ _04717_ _04118_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__nor2_1
XFILLER_6_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17872_ _09684_ _09389_ vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__nand2_1
XFILLER_227_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19611_ rbzero.debug_overlay.playerX\[0\] _02981_ _02985_ _02978_ vssd1 vssd1 vccd1
+ vccd1 _00969_ sky130_fd_sc_hd__o211a_1
XFILLER_120_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16823_ _09364_ _09358_ _09362_ _09363_ vssd1 vssd1 vccd1 vccd1 _09366_ sky130_fd_sc_hd__a211oi_2
XFILLER_24_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19542_ rbzero.pov.spi_buffer\[66\] rbzero.pov.spi_buffer\[67\] _02932_ vssd1 vssd1
+ vccd1 vccd1 _02940_ sky130_fd_sc_hd__mux2_1
XFILLER_219_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13966_ _06648_ _06654_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__nor2_1
XFILLER_171_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16754_ rbzero.wall_tracer.trackDistX\[-9\] rbzero.wall_tracer.stepDistX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _09305_ sky130_fd_sc_hd__nand2_1
XFILLER_235_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15705_ _08271_ _08314_ _08318_ vssd1 vssd1 vccd1 vccd1 _08319_ sky130_fd_sc_hd__nor3_1
X_12917_ _05567_ _05583_ _05605_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__and3_1
XFILLER_34_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16685_ _09257_ vssd1 vssd1 vccd1 vccd1 _09263_ sky130_fd_sc_hd__buf_2
X_19473_ rbzero.pov.spi_buffer\[33\] rbzero.pov.spi_buffer\[34\] _02899_ vssd1 vssd1
+ vccd1 vccd1 _02904_ sky130_fd_sc_hd__mux2_1
XFILLER_234_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13897_ _05434_ _06137_ _06305_ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__or3_1
XFILLER_234_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18424_ _02175_ _02162_ _02161_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a21oi_1
XFILLER_221_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15636_ _08196_ _08206_ vssd1 vssd1 vccd1 vccd1 _08250_ sky130_fd_sc_hd__or2_1
X_12848_ _05527_ _05457_ _05533_ _05536_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__a211oi_4
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18355_ _02107_ _02109_ _02108_ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__o21bai_1
X_15567_ _07378_ _07507_ _07592_ _07399_ vssd1 vssd1 vccd1 vccd1 _08181_ sky130_fd_sc_hd__o22ai_1
XFILLER_37_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12779_ _05460_ _05464_ _05466_ _05467_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__o211a_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17306_ _09828_ _09844_ vssd1 vssd1 vccd1 vccd1 _09845_ sky130_fd_sc_hd__xor2_1
X_14518_ rbzero.wall_tracer.stepDistY\[-2\] _07196_ _07193_ vssd1 vssd1 vccd1 vccd1
+ _07197_ sky130_fd_sc_hd__mux2_1
XFILLER_222_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18286_ _02052_ _02053_ _02054_ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__a21oi_1
X_15498_ _08073_ _08106_ vssd1 vssd1 vccd1 vccd1 _08112_ sky130_fd_sc_hd__xor2_1
XFILLER_175_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17237_ _09652_ _09658_ _09775_ vssd1 vssd1 vccd1 vccd1 _09776_ sky130_fd_sc_hd__o21ai_1
XFILLER_174_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14449_ rbzero.wall_tracer.stepDistY\[-11\] _07136_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _07137_ sky130_fd_sc_hd__mux2_1
XFILLER_70_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17168_ _09577_ _09706_ _09707_ _09576_ vssd1 vssd1 vccd1 vccd1 _09708_ sky130_fd_sc_hd__a22o_1
XFILLER_174_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16119_ _08599_ _08668_ vssd1 vssd1 vccd1 vccd1 _08731_ sky130_fd_sc_hd__or2_1
XFILLER_143_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17099_ _09638_ _09639_ vssd1 vssd1 vccd1 vccd1 _09640_ sky130_fd_sc_hd__xnor2_4
XFILLER_192_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19809_ _02863_ vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__clkinv_2
XFILLER_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20515_ net129 _00531_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20446_ net125 _00477_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20377_ net120 _00408_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13820_ _06467_ _06508_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13751_ _05738_ _06305_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__nand2_1
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10963_ _03709_ vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12702_ _05298_ _05300_ _05307_ _05309_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__nand4_1
XFILLER_147_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16470_ _08903_ _08944_ _09079_ vssd1 vssd1 vccd1 vccd1 _09080_ sky130_fd_sc_hd__a21bo_1
XFILLER_203_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13682_ _06370_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__inv_2
XFILLER_44_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10894_ _03673_ vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15421_ _07961_ _08034_ vssd1 vssd1 vccd1 vccd1 _08035_ sky130_fd_sc_hd__xnor2_2
X_12633_ _05314_ _05318_ _05321_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__and3b_1
XFILLER_223_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18140_ _01919_ _01920_ _09275_ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__o21a_1
XFILLER_180_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15352_ _07416_ _07575_ vssd1 vssd1 vccd1 vccd1 _07966_ sky130_fd_sc_hd__nor2_1
XFILLER_129_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12564_ rbzero.wall_tracer.rayAddendX\[-4\] _05252_ _05219_ vssd1 vssd1 vccd1 vccd1
+ _05253_ sky130_fd_sc_hd__mux2_4
XFILLER_196_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14303_ _06402_ _06982_ vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__xor2_1
XFILLER_54_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18071_ _01732_ _01851_ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__xnor2_1
X_11515_ _04203_ _04207_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__and2_1
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15283_ _07894_ _07895_ vssd1 vssd1 vccd1 vccd1 _07897_ sky130_fd_sc_hd__nand2_1
XFILLER_156_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12495_ _05181_ _05182_ rbzero.debug_overlay.facingX\[10\] _05183_ vssd1 vssd1 vccd1
+ vccd1 _05184_ sky130_fd_sc_hd__a2bb2o_4
X_17022_ _09443_ _09528_ _09562_ vssd1 vssd1 vccd1 vccd1 _09563_ sky130_fd_sc_hd__a21oi_1
X_14234_ _06921_ _06922_ vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__nor2_1
XFILLER_144_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11446_ _04160_ _04163_ _03923_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__mux2_1
XFILLER_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14165_ _06845_ _06848_ _06850_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__nand3_1
XFILLER_67_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11377_ _04067_ _04069_ _04095_ _03295_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13116_ _05766_ _05567_ _05748_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__and3_1
XFILLER_153_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10328_ rbzero.tex_r1\[60\] rbzero.tex_r1\[61\] _03366_ vssd1 vssd1 vccd1 vccd1 _03374_
+ sky130_fd_sc_hd__mux2_1
X_14096_ _06683_ _06681_ vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__xor2_1
X_18973_ _02646_ vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__clkbuf_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17924_ _10155_ _01706_ _01521_ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__o21a_1
X_13047_ _05666_ _05697_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__or2b_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ rbzero.tex_b1\[29\] rbzero.tex_b1\[30\] _03333_ vssd1 vssd1 vccd1 vccd1 _03338_
+ sky130_fd_sc_hd__mux2_1
XTAP_6970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17855_ _01574_ _01636_ _01637_ _09978_ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_121_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16806_ _04940_ vssd1 vssd1 vccd1 vccd1 _09351_ sky130_fd_sc_hd__clkbuf_4
XFILLER_66_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17786_ _01568_ _01569_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__nand2_1
XFILLER_81_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14998_ _07605_ _07611_ vssd1 vssd1 vccd1 vccd1 _07612_ sky130_fd_sc_hd__nand2_1
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19525_ rbzero.pov.spi_buffer\[58\] rbzero.pov.spi_buffer\[59\] _02921_ vssd1 vssd1
+ vccd1 vccd1 _02931_ sky130_fd_sc_hd__mux2_1
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16737_ _09287_ _09288_ _09280_ vssd1 vssd1 vccd1 vccd1 _09290_ sky130_fd_sc_hd__a21bo_1
XFILLER_35_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13949_ _06581_ _06637_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__and2_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19456_ rbzero.pov.spi_buffer\[25\] rbzero.pov.spi_buffer\[26\] _02888_ vssd1 vssd1
+ vccd1 vccd1 _02895_ sky130_fd_sc_hd__mux2_1
X_16668_ rbzero.row_render.size\[5\] _09255_ _07192_ _09259_ vssd1 vssd1 vccd1 vccd1
+ _00503_ sky130_fd_sc_hd__a22o_1
XFILLER_222_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18407_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__nor2_1
X_15619_ _07378_ _07592_ vssd1 vssd1 vccd1 vccd1 _08233_ sky130_fd_sc_hd__or2_1
XFILLER_50_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19387_ _02861_ vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__clkinv_2
X_16599_ _08785_ _09207_ _07835_ vssd1 vssd1 vccd1 vccd1 _09208_ sky130_fd_sc_hd__a21oi_1
XFILLER_188_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18338_ _05001_ _02001_ _02100_ vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__a21oi_1
XFILLER_241_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18269_ rbzero.wall_tracer.trackDistY\[-5\] rbzero.wall_tracer.stepDistY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__nand2_1
XFILLER_50_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20300_ _03258_ vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__clkinv_2
XFILLER_129_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21280_ _00329_ _01296_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20231_ rbzero.traced_texa\[9\] rbzero.texV\[9\] _03242_ vssd1 vssd1 vccd1 vccd1
+ _03247_ sky130_fd_sc_hd__a21o_1
XFILLER_11_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20162_ rbzero.traced_texa\[-1\] rbzero.texV\[-1\] vssd1 vssd1 vccd1 vccd1 _03189_
+ sky130_fd_sc_hd__nand2_1
XFILLER_118_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20093_ gpout5.clk_div\[1\] gpout5.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__nand2_1
XFILLER_170_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20995_ net66 _01011_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_225_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11300_ rbzero.tex_r0\[7\] rbzero.tex_r0\[6\] _03961_ vssd1 vssd1 vccd1 vccd1 _04019_
+ sky130_fd_sc_hd__mux2_1
XFILLER_193_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12280_ rbzero.wall_tracer.trackDistY\[-8\] _04963_ _04965_ rbzero.wall_tracer.trackDistY\[-9\]
+ _04973_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__o221a_1
XFILLER_138_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11231_ _03949_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__clkbuf_4
XFILLER_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20429_ net117 _00460_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11162_ rbzero.traced_texVinit\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _03881_
+ sky130_fd_sc_hd__or2_1
XTAP_6211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15970_ _07343_ _07491_ vssd1 vssd1 vccd1 vccd1 _08584_ sky130_fd_sc_hd__or2_1
X_11093_ _03730_ _03814_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__nor2_1
XFILLER_216_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14921_ _07534_ rbzero.debug_overlay.playerY\[-3\] _05113_ vssd1 vssd1 vccd1 vccd1
+ _07535_ sky130_fd_sc_hd__mux2_1
XTAP_6299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17640_ _10173_ _10174_ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__nand2_1
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14852_ _07356_ vssd1 vssd1 vccd1 vccd1 _07466_ sky130_fd_sc_hd__buf_4
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13803_ _06408_ _06459_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__or2b_1
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17571_ _10093_ _10107_ vssd1 vssd1 vccd1 vccd1 _10108_ sky130_fd_sc_hd__xor2_1
X_14783_ _04935_ _07396_ vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__nand2_1
XFILLER_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11995_ _04694_ _04704_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__nor2_1
XFILLER_216_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19310_ _02840_ _02841_ _02844_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__and3b_1
X_16522_ _08592_ _08296_ _07916_ _08716_ vssd1 vssd1 vccd1 vccd1 _09131_ sky130_fd_sc_hd__or4_1
XFILLER_205_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13734_ _06422_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__clkbuf_4
XFILLER_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10946_ _03700_ vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19241_ rbzero.spi_registers.spi_cmd\[0\] _02784_ rbzero.spi_registers.spi_cmd\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__or3b_1
XFILLER_108_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16453_ _09059_ _09060_ _09062_ vssd1 vssd1 vccd1 vccd1 _09063_ sky130_fd_sc_hd__nand3_1
XFILLER_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13665_ _06348_ _06349_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__xnor2_1
XFILLER_220_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10877_ _03664_ vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _08014_ _08016_ _08017_ vssd1 vssd1 vccd1 vccd1 _08018_ sky130_fd_sc_hd__a21o_1
X_12616_ _05296_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__clkbuf_4
X_16384_ _08982_ _08993_ vssd1 vssd1 vccd1 vccd1 _08994_ sky130_fd_sc_hd__xor2_1
XFILLER_188_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19172_ _09247_ _02761_ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__and2_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _06263_ _06284_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__and2_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18123_ _01901_ _01903_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__or2_1
X_15335_ _07933_ _07946_ vssd1 vssd1 vccd1 vccd1 _07949_ sky130_fd_sc_hd__nor2_1
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12547_ _05234_ _05235_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__xnor2_2
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18054_ _01733_ _01753_ _01731_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__a21o_1
X_15266_ _07879_ vssd1 vssd1 vccd1 vccd1 _07880_ sky130_fd_sc_hd__clkbuf_4
XFILLER_145_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12478_ _05165_ _05166_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__and2b_1
XANTENNA_3 _02720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17005_ _09408_ _09410_ _09407_ vssd1 vssd1 vccd1 vccd1 _09546_ sky130_fd_sc_hd__a21bo_1
XFILLER_201_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14217_ _06885_ _06905_ vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__nand2_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11429_ _03968_ _04140_ _04141_ _04146_ _03972_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__o221a_1
X_15197_ _07787_ _07810_ vssd1 vssd1 vccd1 vccd1 _07811_ sky130_fd_sc_hd__xor2_1
XFILLER_119_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14148_ _06796_ _06797_ _06834_ vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__a21o_1
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14079_ _06766_ _06767_ vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__xnor2_1
X_18956_ _02637_ vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__clkbuf_1
XFILLER_234_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17907_ _01688_ _01689_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__nor2_1
XFILLER_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18887_ _02590_ _02597_ _02598_ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__and3_1
XFILLER_230_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17838_ _01588_ _01620_ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__xor2_2
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17769_ _09829_ _08735_ vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__nor2_1
XFILLER_78_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19508_ _02922_ vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20780_ net87 _00796_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19439_ rbzero.pov.spi_buffer\[17\] rbzero.pov.spi_buffer\[18\] _02877_ vssd1 vssd1
+ vccd1 vccd1 _02886_ sky130_fd_sc_hd__mux2_1
XFILLER_223_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21401_ net86 _01417_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_202_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21332_ _00355_ _01348_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21263_ _00312_ _01279_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20214_ _03231_ _03232_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21194_ _00243_ _01210_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20145_ rbzero.traced_texa\[-5\] rbzero.texV\[-5\] _03174_ vssd1 vssd1 vccd1 vccd1
+ _03175_ sky130_fd_sc_hd__o21ai_1
XFILLER_213_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ _03130_ vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__clkinv_2
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ rbzero.tex_g0\[31\] rbzero.tex_g0\[30\] _03616_ vssd1 vssd1 vccd1 vccd1 _03624_
+ sky130_fd_sc_hd__mux2_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ rbzero.tex_b0\[23\] _04143_ _04145_ _03930_ vssd1 vssd1 vccd1 vccd1 _04495_
+ sky130_fd_sc_hd__a31o_1
XFILLER_57_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20978_ net64 _00994_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10731_ _03587_ vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13450_ _06133_ _06131_ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__nor2_1
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10662_ _03551_ vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12401_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__nand2_1
XFILLER_224_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13381_ _06069_ _06051_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10593_ _03515_ vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15120_ _04935_ rbzero.wall_tracer.stepDistX\[-2\] vssd1 vssd1 vccd1 vccd1 _07734_
+ sky130_fd_sc_hd__nand2_1
XFILLER_154_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12332_ _03801_ _03779_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__and2_2
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15051_ _07663_ _07664_ vssd1 vssd1 vccd1 vccd1 _07665_ sky130_fd_sc_hd__nor2_1
X_12263_ _04945_ rbzero.wall_tracer.trackDistX\[0\] vssd1 vssd1 vccd1 vccd1 _04957_
+ sky130_fd_sc_hd__and2_1
XFILLER_120_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14002_ _06137_ _06343_ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__nor2_1
XFILLER_107_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11214_ rbzero.tex_r0\[57\] rbzero.tex_r0\[56\] _03925_ vssd1 vssd1 vccd1 vccd1 _03933_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12194_ net34 _04874_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__and2b_1
XFILLER_107_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18810_ _02507_ _02508_ _02517_ vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__nor3_1
XTAP_6030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11145_ _03852_ _03860_ _03863_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__o21a_1
XTAP_6041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19790_ _03085_ _03091_ _03092_ _03093_ _04101_ vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__a32o_1
XFILLER_7_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18741_ _02440_ _02450_ vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__nand2_1
XTAP_6085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11076_ _03799_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__clkbuf_4
XTAP_5340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15953_ _08565_ _08566_ vssd1 vssd1 vccd1 vccd1 _08567_ sky130_fd_sc_hd__nand2_1
XFILLER_7_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14904_ _07501_ _07508_ _07510_ _07517_ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__or4_1
XTAP_5373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18672_ _02401_ _02389_ _02387_ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__a21oi_1
XFILLER_248_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15884_ _08471_ _08496_ _08497_ vssd1 vssd1 vccd1 vccd1 _08498_ sky130_fd_sc_hd__nand3_1
XTAP_5395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17623_ _10087_ _10153_ _10157_ vssd1 vssd1 vccd1 vccd1 _10159_ sky130_fd_sc_hd__and3_1
X_14835_ _07446_ _07447_ _07448_ vssd1 vssd1 vccd1 vccd1 _07449_ sky130_fd_sc_hd__or3_1
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _09967_ _09969_ vssd1 vssd1 vccd1 vccd1 _10091_ sky130_fd_sc_hd__nor2_1
XFILLER_189_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14766_ _07355_ _07379_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__nor2_1
X_11978_ net19 _04686_ _04687_ net18 vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__a31o_1
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16505_ _09113_ vssd1 vssd1 vccd1 vccd1 _09114_ sky130_fd_sc_hd__buf_2
X_13717_ _05641_ _06304_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__and2_1
X_10929_ _03691_ vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__clkbuf_1
X_17485_ _09369_ _09761_ _10022_ vssd1 vssd1 vccd1 vccd1 _10023_ sky130_fd_sc_hd__a21o_1
X_14697_ rbzero.wall_tracer.stepDistX\[3\] _07211_ _07316_ vssd1 vssd1 vccd1 vccd1
+ _07323_ sky130_fd_sc_hd__mux2_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19224_ rbzero.spi_registers.got_new_sky _02742_ _02740_ _02793_ vssd1 vssd1 vccd1
+ vccd1 _00774_ sky130_fd_sc_hd__a31o_1
X_16436_ _09035_ _09045_ vssd1 vssd1 vccd1 vccd1 _09046_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13648_ _06306_ _06335_ _06336_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__and3_1
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19155_ rbzero.spi_registers.new_leak\[5\] _02745_ vssd1 vssd1 vccd1 vccd1 _02751_
+ sky130_fd_sc_hd__or2_1
X_16367_ _08902_ _08883_ vssd1 vssd1 vccd1 vccd1 _08977_ sky130_fd_sc_hd__or2b_1
X_13579_ _05645_ _05701_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__nand2_1
XFILLER_121_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18106_ _01856_ _01886_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__xnor2_1
XFILLER_160_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15318_ _07773_ _07779_ vssd1 vssd1 vccd1 vccd1 _07932_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16298_ _08907_ _08908_ vssd1 vssd1 vccd1 vccd1 _08909_ sky130_fd_sc_hd__xnor2_1
X_19086_ _02706_ vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18037_ _01728_ _01729_ _01817_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__and3_1
X_15249_ _07379_ _07712_ _07736_ _07400_ vssd1 vssd1 vccd1 vccd1 _07863_ sky130_fd_sc_hd__o22a_1
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19988_ _03121_ vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__clkinv_2
XFILLER_98_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18939_ _02628_ vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__clkbuf_1
XFILLER_234_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20901_ net60 _00917_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20832_ _00050_ _00848_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20763_ net107 _00779_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20694_ net84 _00710_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_167_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21315_ _00338_ _01331_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21246_ _00295_ _01262_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21177_ _00226_ _01193_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_77_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20128_ _03158_ _03159_ _03160_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__nand3_1
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12950_ _05608_ _05638_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__nor2_1
XFILLER_218_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20059_ _03125_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__buf_4
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11901_ _04611_ o_rgb[14] vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__or2_1
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _05531_ _05504_ _05569_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__o21a_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _07275_ _07254_ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__nor2_1
X_11832_ rbzero.tex_b1\[37\] rbzero.tex_b1\[36\] _04032_ vssd1 vssd1 vccd1 vccd1 _04546_
+ sky130_fd_sc_hd__mux2_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14551_ _07222_ vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__clkbuf_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11763_ _03957_ _04475_ _04476_ _04477_ _03946_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__o221a_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13502_ _06182_ _06190_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__nand2_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ rbzero.tex_g1\[7\] rbzero.tex_g1\[8\] _03574_ vssd1 vssd1 vccd1 vccd1 _03579_
+ sky130_fd_sc_hd__mux2_1
X_17270_ _09702_ _09704_ _09701_ vssd1 vssd1 vccd1 vccd1 _09809_ sky130_fd_sc_hd__a21oi_1
X_14482_ _07166_ vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__clkbuf_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11694_ rbzero.tex_g1\[63\] rbzero.tex_g1\[62\] _04378_ vssd1 vssd1 vccd1 vccd1 _04410_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13433_ _05612_ _05525_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__xnor2_1
X_16221_ _08831_ _08832_ vssd1 vssd1 vccd1 vccd1 _08833_ sky130_fd_sc_hd__nor2_1
XFILLER_201_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10645_ rbzero.tex_g1\[40\] rbzero.tex_g1\[41\] _03541_ vssd1 vssd1 vccd1 vccd1 _03543_
+ sky130_fd_sc_hd__mux2_1
XFILLER_195_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16152_ _08748_ _08624_ _08763_ vssd1 vssd1 vccd1 vccd1 _08764_ sky130_fd_sc_hd__a21o_1
XFILLER_195_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13364_ _06049_ _06051_ _06052_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__a21oi_1
XFILLER_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10576_ _03506_ vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__clkbuf_1
X_12315_ _05001_ rbzero.wall_tracer.trackDistX\[4\] _05006_ _05007_ _05008_ vssd1
+ vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__a2111o_1
X_15103_ _07709_ _07710_ _07646_ vssd1 vssd1 vccd1 vccd1 _07717_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16083_ _08693_ _08695_ vssd1 vssd1 vccd1 vccd1 _08696_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13295_ _05615_ _05982_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__xnor2_1
XFILLER_182_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15034_ _07208_ _07445_ vssd1 vssd1 vccd1 vccd1 _07648_ sky130_fd_sc_hd__xnor2_4
XFILLER_177_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19911_ _03113_ vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__clkinv_2
X_12246_ _03731_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__buf_6
XFILLER_29_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19842_ _03107_ vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__clkinv_2
X_12177_ _04874_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__buf_2
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ _03844_ _03843_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__nand2_1
X_19773_ _03289_ _03443_ _03080_ _03078_ _04920_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__o41a_1
XFILLER_231_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16985_ _09376_ _09525_ vssd1 vssd1 vccd1 vccd1 _09526_ sky130_fd_sc_hd__xor2_1
XFILLER_49_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18724_ _02448_ _02449_ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__nand2_1
X_15936_ _08548_ _08549_ vssd1 vssd1 vccd1 vccd1 _08550_ sky130_fd_sc_hd__nand2_1
XTAP_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11059_ _03291_ _03294_ _03296_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__or3_1
XFILLER_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18655_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.wall_tracer.rayAddendY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__nor2_1
X_15867_ _08472_ _08479_ _08480_ vssd1 vssd1 vccd1 vccd1 _08481_ sky130_fd_sc_hd__and3_1
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17606_ _10036_ _10037_ _10142_ vssd1 vssd1 vccd1 vccd1 _10143_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14818_ rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18586_ rbzero.wall_tracer.rayAddendX\[8\] rbzero.wall_tracer.rayAddendX\[7\] _02275_
+ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__o21a_1
X_15798_ _08323_ _08350_ vssd1 vssd1 vccd1 vccd1 _08412_ sky130_fd_sc_hd__nand2_1
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_152 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_152/HI o_rgb[12]
+ sky130_fd_sc_hd__conb_1
XFILLER_205_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17537_ _08732_ _09829_ vssd1 vssd1 vccd1 vccd1 _10074_ sky130_fd_sc_hd__nor2_1
X_14749_ rbzero.wall_tracer.visualWallDist\[-6\] _03793_ vssd1 vssd1 vccd1 vccd1 _07363_
+ sky130_fd_sc_hd__and2_1
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17468_ _09870_ _09872_ vssd1 vssd1 vccd1 vccd1 _10006_ sky130_fd_sc_hd__nor2_1
XFILLER_178_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19207_ _02783_ vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16419_ _09027_ _09028_ vssd1 vssd1 vccd1 vccd1 _09029_ sky130_fd_sc_hd__xor2_1
XFILLER_220_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17399_ _09935_ _09936_ vssd1 vssd1 vccd1 vccd1 _09937_ sky130_fd_sc_hd__nand2_1
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19138_ _04111_ _04252_ _04113_ _02719_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__nand4_4
XFILLER_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19069_ rbzero.spi_registers.spi_buffer\[6\] rbzero.spi_registers.spi_buffer\[5\]
+ _02690_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__mux2_1
XFILLER_218_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21100_ _00149_ _01116_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21031_ net101 _01047_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_vinf
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout104 net108 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__buf_2
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout115 net141 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_4
XFILLER_232_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout126 net141 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout137 net139 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_2
XFILLER_247_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20815_ _00033_ _00831_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20746_ net103 _00762_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20677_ net67 _00693_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10430_ rbzero.tex_r1\[12\] rbzero.tex_r1\[13\] _03422_ vssd1 vssd1 vccd1 vccd1 _03428_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10361_ rbzero.tex_r1\[45\] rbzero.tex_r1\[46\] _03389_ vssd1 vssd1 vccd1 vccd1 _03392_
+ sky130_fd_sc_hd__mux2_1
XFILLER_104_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12100_ _04785_ net23 _04801_ _04807_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__a31o_1
XFILLER_30_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13080_ _05766_ _05722_ _05768_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__and3_1
XFILLER_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10292_ _03299_ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12031_ _03784_ _03291_ gpout0.vpos\[6\] gpout0.vpos\[7\] net3 _04731_ vssd1 vssd1
+ vccd1 vccd1 _04740_ sky130_fd_sc_hd__mux4_1
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21229_ _00278_ _01245_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16770_ rbzero.wall_tracer.trackDistX\[-7\] rbzero.wall_tracer.stepDistX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _09319_ sky130_fd_sc_hd__nand2_1
XFILLER_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13982_ _06516_ _06668_ _06670_ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__a21bo_1
XFILLER_120_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15721_ _07718_ vssd1 vssd1 vccd1 vccd1 _08335_ sky130_fd_sc_hd__buf_4
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ _05526_ _05545_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__xnor2_4
XFILLER_20_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ rbzero.debug_overlay.vplaneX\[-1\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__or2_1
X_15652_ _08249_ _08250_ _08262_ _08263_ _08265_ vssd1 vssd1 vccd1 vccd1 _08266_ sky130_fd_sc_hd__a32o_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _05552_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__clkinv_2
XFILLER_2_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _05016_ _07254_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__nor2_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _02125_ _02126_ _02127_ _09351_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__a31o_1
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11815_ _04527_ _04528_ _03928_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__mux2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _08135_ _08136_ vssd1 vssd1 vccd1 vccd1 _08197_ sky130_fd_sc_hd__nand2_1
X_12795_ _05422_ _05450_ _05448_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__mux2_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _09476_ _09609_ _09732_ _09734_ vssd1 vssd1 vccd1 vccd1 _09861_ sky130_fd_sc_hd__and4b_2
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14534_ rbzero.wall_tracer.stepDistY\[2\] _07208_ _07193_ vssd1 vssd1 vccd1 vccd1
+ _07209_ sky130_fd_sc_hd__mux2_1
X_11746_ rbzero.tex_b0\[53\] rbzero.tex_b0\[52\] _03959_ vssd1 vssd1 vccd1 vccd1 _04461_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17253_ _08596_ _08851_ _09373_ _08599_ vssd1 vssd1 vccd1 vccd1 _09792_ sky130_fd_sc_hd__o22a_1
XFILLER_202_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14465_ _07127_ _07120_ _07105_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__mux2_1
X_11677_ rbzero.tex_g1\[2\] _04374_ _03997_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__a21o_1
XFILLER_169_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16204_ _08658_ _08685_ _08815_ vssd1 vssd1 vccd1 vccd1 _08816_ sky130_fd_sc_hd__a21oi_1
XFILLER_179_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13416_ _06028_ _05738_ _06102_ _06103_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__a22o_1
XFILLER_128_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10628_ rbzero.tex_g1\[48\] rbzero.tex_g1\[49\] _03530_ vssd1 vssd1 vccd1 vccd1 _03534_
+ sky130_fd_sc_hd__mux2_1
X_17184_ _07858_ _09451_ vssd1 vssd1 vccd1 vccd1 _09724_ sky130_fd_sc_hd__nor2_1
X_14396_ _07067_ _07084_ _05531_ vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__mux2_1
XFILLER_174_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16135_ _08601_ _08610_ _08609_ vssd1 vssd1 vccd1 vccd1 _08747_ sky130_fd_sc_hd__a21o_1
X_13347_ _06030_ _06031_ _06035_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10559_ _03497_ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16066_ _08677_ _08678_ vssd1 vssd1 vccd1 vccd1 _08679_ sky130_fd_sc_hd__nor2_1
XFILLER_192_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13278_ _05962_ _05965_ _05966_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__and3_1
XFILLER_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15017_ _07524_ vssd1 vssd1 vccd1 vccd1 _07631_ sky130_fd_sc_hd__clkbuf_4
XFILLER_170_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12229_ _04926_ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19825_ _03105_ vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__clkinv_2
XFILLER_25_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19756_ rbzero.pov.ready_buffer\[6\] _03067_ _03068_ rbzero.debug_overlay.vplaneY\[-3\]
+ _03015_ vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__a221o_1
X_16968_ rbzero.wall_tracer.trackDistX\[0\] rbzero.wall_tracer.stepDistX\[0\] vssd1
+ vssd1 vccd1 vccd1 _09510_ sky130_fd_sc_hd__nand2_1
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18707_ _02414_ _02424_ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__nand2_1
XFILLER_204_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15919_ _07913_ _07917_ _07911_ vssd1 vssd1 vccd1 vccd1 _08533_ sky130_fd_sc_hd__a21o_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19687_ _03043_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__inv_2
XFILLER_83_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16899_ _09438_ _09440_ vssd1 vssd1 vccd1 vccd1 _09441_ sky130_fd_sc_hd__xor2_1
X_18638_ _02370_ vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18569_ _02309_ _02310_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__nand2_1
XFILLER_52_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20600_ net82 _00616_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_205_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20531_ net121 _00547_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20462_ net96 _00478_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.wall\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20393_ net138 _00424_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_161_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21014_ net81 _01030_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11600_ _03972_ _04312_ _04316_ _03950_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__a211o_1
XFILLER_70_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12580_ rbzero.wall_tracer.visualWallDist\[0\] _05190_ _03789_ vssd1 vssd1 vccd1
+ vccd1 _05269_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11531_ rbzero.debug_overlay.facingX\[-9\] _04240_ _04242_ rbzero.debug_overlay.facingX\[-4\]
+ _04248_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__a221o_1
XFILLER_8_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20729_ net100 _00745_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14250_ _06935_ _06936_ _06938_ vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__o21a_1
XFILLER_8_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11462_ rbzero.tex_r1\[10\] _03961_ _03929_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__a21o_1
XFILLER_165_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13201_ _05692_ _05641_ _05886_ _05889_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__a31o_1
XFILLER_104_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10413_ rbzero.tex_r1\[20\] rbzero.tex_r1\[21\] _03411_ vssd1 vssd1 vccd1 vccd1 _03419_
+ sky130_fd_sc_hd__mux2_1
X_14181_ _06868_ _06869_ vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__and2b_1
XFILLER_183_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11393_ gpout0.vpos\[8\] gpout0.vpos\[7\] gpout0.vpos\[6\] vssd1 vssd1 vccd1 vccd1
+ _04112_ sky130_fd_sc_hd__and3_1
XFILLER_125_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13132_ _05671_ _05728_ _05726_ _05629_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__o22a_1
X_10344_ _03382_ vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17940_ rbzero.wall_tracer.trackDistX\[8\] rbzero.wall_tracer.stepDistX\[8\] vssd1
+ vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__nand2_1
X_13063_ _05608_ _05611_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__nor2_1
XFILLER_112_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10275_ _03346_ vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_239_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12014_ _04717_ o_rgb[14] _04722_ net7 vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__o211a_1
XFILLER_79_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17871_ _01652_ _01653_ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__or2b_1
XFILLER_117_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19610_ rbzero.pov.ready_buffer\[68\] _02836_ _02955_ _02984_ vssd1 vssd1 vccd1 vccd1
+ _02985_ sky130_fd_sc_hd__a211o_1
X_16822_ _09362_ _09363_ _09364_ _09358_ vssd1 vssd1 vccd1 vccd1 _09365_ sky130_fd_sc_hd__o211a_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19541_ _02939_ vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__clkbuf_1
XFILLER_235_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16753_ rbzero.wall_tracer.trackDistX\[-9\] rbzero.wall_tracer.stepDistX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _09304_ sky130_fd_sc_hd__or2_1
XFILLER_24_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13965_ _06596_ _06649_ _06650_ _06653_ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_150_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15704_ _08315_ _08317_ vssd1 vssd1 vccd1 vccd1 _08318_ sky130_fd_sc_hd__xnor2_2
XFILLER_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12916_ _05591_ _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__nor2_1
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19472_ _02903_ vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__clkbuf_1
X_16684_ rbzero.traced_texa\[-11\] _09262_ _09258_ rbzero.wall_tracer.visualWallDist\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__a22o_1
XFILLER_98_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13896_ _06547_ _06584_ vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__or2_1
XFILLER_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18423_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__or2_1
XFILLER_234_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15635_ _08196_ _08206_ vssd1 vssd1 vccd1 vccd1 _08249_ sky130_fd_sc_hd__nand2_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12847_ _05499_ _05465_ _05534_ _05535_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__o211a_1
XFILLER_37_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18354_ rbzero.wall_tracer.trackDistY\[7\] rbzero.wall_tracer.stepDistY\[7\] vssd1
+ vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__nand2_1
XFILLER_199_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15566_ _07416_ _07986_ vssd1 vssd1 vccd1 vccd1 _08180_ sky130_fd_sc_hd__nor2_1
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12778_ _05404_ _05445_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__nand2_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _09835_ _09843_ vssd1 vssd1 vccd1 vccd1 _09844_ sky130_fd_sc_hd__xnor2_1
XFILLER_226_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14517_ _07102_ _07195_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__nand2_1
X_18285_ _02052_ _02053_ _02054_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__and3_1
X_11729_ rbzero.color_sky\[3\] rbzero.color_floor\[3\] _04030_ vssd1 vssd1 vccd1 vccd1
+ _04445_ sky130_fd_sc_hd__mux2_1
XFILLER_222_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15497_ _08036_ _08108_ vssd1 vssd1 vccd1 vccd1 _08111_ sky130_fd_sc_hd__xor2_1
X_17236_ _09520_ _09659_ vssd1 vssd1 vccd1 vccd1 _09775_ sky130_fd_sc_hd__nand2_1
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14448_ _07102_ _07135_ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__nand2_1
XFILLER_204_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17167_ _07824_ _08793_ _07890_ vssd1 vssd1 vccd1 vccd1 _09707_ sky130_fd_sc_hd__a21o_1
X_14379_ _07029_ _07067_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__nor2_1
XFILLER_128_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16118_ _08597_ _08600_ _08593_ vssd1 vssd1 vccd1 vccd1 _08730_ sky130_fd_sc_hd__a21bo_1
XFILLER_157_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17098_ _09369_ _09506_ _09504_ vssd1 vssd1 vccd1 vccd1 _09639_ sky130_fd_sc_hd__a21oi_2
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16049_ _08429_ _08531_ vssd1 vssd1 vccd1 vccd1 _08662_ sky130_fd_sc_hd__or2_1
XFILLER_192_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19808_ rbzero.spi_registers.got_new_vinf _02742_ _02740_ _02141_ vssd1 vssd1 vccd1
+ vccd1 _01047_ sky130_fd_sc_hd__a31o_1
XFILLER_245_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19739_ rbzero.pov.ready_buffer\[11\] _03069_ _03070_ rbzero.debug_overlay.vplaneX\[-9\]
+ _03065_ vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__o221a_1
XFILLER_237_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20514_ net129 _00530_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20445_ net139 _00476_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20376_ net124 _00407_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_161_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_7127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13750_ _06410_ _06415_ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10962_ rbzero.tex_b0\[18\] rbzero.tex_b0\[17\] _03704_ vssd1 vssd1 vccd1 vccd1 _03709_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12701_ _05351_ _05354_ _05389_ _05387_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__or4_1
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13681_ _06367_ _06369_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__and2b_1
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10893_ rbzero.tex_b0\[51\] rbzero.tex_b0\[50\] _03671_ vssd1 vssd1 vccd1 vccd1 _03673_
+ sky130_fd_sc_hd__mux2_1
XFILLER_231_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15420_ _08002_ _08032_ _08033_ vssd1 vssd1 vccd1 vccd1 _08034_ sky130_fd_sc_hd__a21oi_2
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12632_ _05319_ _05320_ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__xnor2_2
XFILLER_231_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15351_ _07378_ _07423_ _07554_ _07964_ vssd1 vssd1 vccd1 vccd1 _07965_ sky130_fd_sc_hd__a2bb2o_1
X_12563_ rbzero.wall_tracer.visualWallDist\[-12\] rbzero.wall_tracer.rayAddendY\[-4\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__mux2_1
XFILLER_145_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14302_ _06986_ _06989_ _06990_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__a21o_1
XFILLER_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11514_ _03780_ _04200_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__and2b_1
X_18070_ _01849_ _01850_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__nor2_1
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15282_ _07894_ _07895_ vssd1 vssd1 vccd1 vccd1 _07896_ sky130_fd_sc_hd__nor2_1
XFILLER_141_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12494_ rbzero.wall_tracer.rayAddendX\[10\] rbzero.wall_tracer.rayAddendX\[9\] vssd1
+ vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__or2_1
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17021_ _09545_ _09561_ vssd1 vssd1 vccd1 vccd1 _09562_ sky130_fd_sc_hd__xnor2_1
X_14233_ _05740_ _06634_ _06389_ _06137_ vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__o22a_1
XFILLER_123_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11445_ _04161_ _04162_ _03910_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__mux2_1
XFILLER_171_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14164_ _06831_ _06852_ vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__or2_1
XFILLER_193_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11376_ _03293_ _04071_ _04073_ _04094_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__o22a_1
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13115_ _05618_ _05745_ _05537_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__a21o_1
X_10327_ _03373_ vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__clkbuf_1
X_14095_ _06706_ _06732_ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__nand2_1
XFILLER_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18972_ rbzero.pov.spi_buffer\[34\] rbzero.pov.ready_buffer\[34\] _02640_ vssd1 vssd1
+ vccd1 vccd1 _02646_ sky130_fd_sc_hd__mux2_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ _01523_ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__inv_2
X_13046_ _05719_ _05734_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__xnor2_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ _03337_ vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17854_ _08241_ _01636_ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__or2_1
XFILLER_67_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10189_ _03301_ vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__clkbuf_1
XFILLER_227_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16805_ _09346_ _09347_ _09348_ vssd1 vssd1 vccd1 vccd1 _09350_ sky130_fd_sc_hd__a21oi_1
X_17785_ _08595_ _08645_ _09055_ _09163_ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14997_ _07607_ _07610_ vssd1 vssd1 vccd1 vccd1 _07611_ sky130_fd_sc_hd__nor2_1
XFILLER_219_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19524_ _02930_ vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16736_ _09280_ _09287_ _09288_ vssd1 vssd1 vccd1 vccd1 _09289_ sky130_fd_sc_hd__nand3b_1
XFILLER_228_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13948_ _05861_ _06634_ _06580_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__o21ai_1
XFILLER_130_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19455_ _02894_ vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__clkbuf_1
X_16667_ rbzero.row_render.size\[4\] _09255_ _07189_ _09259_ vssd1 vssd1 vccd1 vccd1
+ _00502_ sky130_fd_sc_hd__a22o_1
XFILLER_234_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13879_ _06564_ _06566_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__nor2_1
XFILLER_50_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18406_ _09258_ _02156_ _02159_ vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__a21o_1
X_15618_ _07416_ _08059_ vssd1 vssd1 vccd1 vccd1 _08232_ sky130_fd_sc_hd__nor2_1
XFILLER_50_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19386_ _02861_ vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__clkinv_2
X_16598_ _04938_ rbzero.wall_tracer.stepDistX\[8\] vssd1 vssd1 vccd1 vccd1 _09207_
+ sky130_fd_sc_hd__nand2_4
XFILLER_210_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18337_ _09351_ _02098_ _02099_ _10028_ _01995_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__o311a_1
X_15549_ _08151_ _08150_ vssd1 vssd1 vccd1 vccd1 _08163_ sky130_fd_sc_hd__and2b_1
XFILLER_163_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18268_ rbzero.wall_tracer.trackDistY\[-5\] rbzero.wall_tracer.stepDistY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__or2_1
XFILLER_200_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17219_ _09758_ vssd1 vssd1 vccd1 vccd1 _09759_ sky130_fd_sc_hd__inv_2
XFILLER_190_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18199_ _01805_ _01977_ _01978_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__o21a_1
XFILLER_116_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20230_ rbzero.traced_texa\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _03246_
+ sky130_fd_sc_hd__nand2_1
XFILLER_144_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20161_ rbzero.traced_texa\[-1\] rbzero.texV\[-1\] vssd1 vssd1 vccd1 vccd1 _03188_
+ sky130_fd_sc_hd__or2_1
XFILLER_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20092_ gpout5.clk_div\[0\] _03003_ vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__nor2_1
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20994_ net56 _01010_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11230_ _03948_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__clkbuf_4
X_20428_ net118 _00459_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11161_ rbzero.traced_texVinit\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _03880_
+ sky130_fd_sc_hd__nand2_1
XFILLER_136_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20359_ gpout3.clk_div\[1\] gpout3.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__nand2_1
XFILLER_84_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11092_ rbzero.wall_tracer.state\[14\] _03813_ rbzero.wall_tracer.state\[10\] vssd1
+ vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__a21oi_1
XTAP_5511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14920_ _07497_ _07533_ vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__and2_1
XTAP_6289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14851_ _07462_ _07464_ _07374_ vssd1 vssd1 vccd1 vccd1 _07465_ sky130_fd_sc_hd__mux2_1
XFILLER_76_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13802_ _06433_ _06490_ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__or2_1
XFILLER_63_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17570_ _10099_ _10106_ vssd1 vssd1 vccd1 vccd1 _10107_ sky130_fd_sc_hd__xnor2_1
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14782_ _07394_ _07395_ _07374_ vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__mux2_1
XFILLER_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11994_ net45 _04697_ _04698_ _04702_ _04703_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__a221o_1
XFILLER_216_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16521_ _08592_ _07916_ _08717_ _08296_ vssd1 vssd1 vccd1 vccd1 _09130_ sky130_fd_sc_hd__o22a_1
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13733_ _06175_ _06421_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__nand2_2
X_10945_ rbzero.tex_b0\[26\] rbzero.tex_b0\[25\] _03693_ vssd1 vssd1 vccd1 vccd1 _03700_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19240_ rbzero.spi_registers.got_new_floor _02742_ _02740_ _02802_ vssd1 vssd1 vccd1
+ vccd1 _00781_ sky130_fd_sc_hd__a31o_1
X_16452_ _07847_ _08787_ _08931_ _09061_ vssd1 vssd1 vccd1 vccd1 _09062_ sky130_fd_sc_hd__o31ai_1
XFILLER_204_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13664_ _05401_ _06352_ _06316_ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__a21o_1
XFILLER_177_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10876_ rbzero.tex_b0\[59\] rbzero.tex_b0\[58\] _03660_ vssd1 vssd1 vccd1 vccd1 _03664_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15403_ _08007_ _08013_ vssd1 vssd1 vccd1 vccd1 _08017_ sky130_fd_sc_hd__nor2_1
XFILLER_231_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ _03790_ _05291_ _05192_ _05187_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__o211ai_1
X_19171_ rbzero.spi_registers.new_sky\[5\] rbzero.color_sky\[5\] _02752_ vssd1 vssd1
+ vccd1 vccd1 _02761_ sky130_fd_sc_hd__mux2_1
XFILLER_231_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16383_ _08991_ _08992_ vssd1 vssd1 vccd1 vccd1 _08993_ sky130_fd_sc_hd__nor2_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13595_ _06265_ _06283_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18122_ _01801_ _01811_ _01902_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__a21oi_1
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15334_ _07488_ _07489_ vssd1 vssd1 vccd1 vccd1 _07948_ sky130_fd_sc_hd__xor2_1
XFILLER_40_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12546_ _05147_ _05154_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__or2b_1
XFILLER_184_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18053_ _01713_ _01716_ _01717_ _01830_ _01833_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__a41o_1
XFILLER_185_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15265_ _07571_ _07572_ vssd1 vssd1 vccd1 vccd1 _07879_ sky130_fd_sc_hd__and2_1
XFILLER_177_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12477_ rbzero.debug_overlay.facingX\[-4\] rbzero.wall_tracer.rayAddendX\[4\] vssd1
+ vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__nand2_1
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17004_ _09535_ _09544_ vssd1 vssd1 vccd1 vccd1 _09545_ sky130_fd_sc_hd__xor2_1
XANTENNA_4 _04026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _06903_ _06904_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__or2_1
XFILLER_172_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11428_ rbzero.tex_r1\[41\] _04143_ _04145_ _03910_ vssd1 vssd1 vccd1 vccd1 _04146_
+ sky130_fd_sc_hd__a31o_1
X_15196_ _07798_ _07809_ vssd1 vssd1 vccd1 vccd1 _07810_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14147_ _06835_ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__inv_2
XFILLER_154_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11359_ gpout0.hpos\[4\] vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__clkbuf_4
XFILLER_119_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14078_ _06101_ _06389_ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__nor2_1
X_18955_ rbzero.pov.spi_buffer\[26\] rbzero.pov.ready_buffer\[26\] _02629_ vssd1 vssd1
+ vccd1 vccd1 _02637_ sky130_fd_sc_hd__mux2_1
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17906_ _01685_ _01687_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__and2_1
X_13029_ _05713_ _05717_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__xnor2_2
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18886_ rbzero.spi_registers.spi_counter\[3\] _02594_ vssd1 vssd1 vccd1 vccd1 _02598_
+ sky130_fd_sc_hd__or2_1
XTAP_6790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17837_ _09182_ _01586_ _01472_ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__o21ai_2
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17768_ _01550_ _01551_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__nand2_1
XFILLER_214_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16719_ _05026_ _09272_ vssd1 vssd1 vccd1 vccd1 _09273_ sky130_fd_sc_hd__and2_1
X_19507_ rbzero.pov.spi_buffer\[49\] rbzero.pov.spi_buffer\[50\] _02921_ vssd1 vssd1
+ vccd1 vccd1 _02922_ sky130_fd_sc_hd__mux2_1
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17699_ _01482_ _01483_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__nor2_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19438_ _02885_ vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19369_ _02859_ vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__clkinv_2
XFILLER_241_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21400_ net86 _01416_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21331_ _00354_ _01347_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21262_ _00311_ _01278_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20213_ _03226_ _03229_ _03227_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21193_ _00242_ _01209_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20144_ rbzero.traced_texa\[-5\] rbzero.texV\[-5\] _03169_ vssd1 vssd1 vccd1 vccd1
+ _03174_ sky130_fd_sc_hd__a21o_1
XFILLER_132_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20075_ _03130_ vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__clkinv_2
XFILLER_246_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20977_ net63 _00993_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10730_ net49 rbzero.tex_g0\[63\] _03512_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__mux2_1
XFILLER_214_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10661_ rbzero.tex_g1\[32\] rbzero.tex_g1\[33\] _03541_ vssd1 vssd1 vccd1 vccd1 _03551_
+ sky130_fd_sc_hd__mux2_1
XFILLER_224_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12400_ _05092_ _05041_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__xnor2_2
XFILLER_22_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13380_ _06048_ _06047_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__xor2_1
X_10592_ rbzero.tex_r0\[2\] rbzero.tex_r0\[1\] _03512_ vssd1 vssd1 vccd1 vccd1 _03515_
+ sky130_fd_sc_hd__mux2_1
XFILLER_222_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ _05011_ _05015_ _05024_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__o21ai_4
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12262_ rbzero.wall_tracer.trackDistX\[-1\] _04953_ vssd1 vssd1 vccd1 vccd1 _04956_
+ sky130_fd_sc_hd__and2_1
X_15050_ rbzero.wall_tracer.visualWallDist\[-11\] _03793_ vssd1 vssd1 vccd1 vccd1
+ _07664_ sky130_fd_sc_hd__nand2_4
XFILLER_108_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14001_ _06631_ _06689_ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11213_ _03909_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__clkbuf_4
XFILLER_108_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12193_ net33 net34 vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__and2b_1
XFILLER_190_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11144_ _03862_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__inv_2
XFILLER_96_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18740_ _02463_ _02464_ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__nor2_1
XFILLER_95_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11075_ _03798_ _03778_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__nand2_2
X_15952_ _08564_ _07344_ vssd1 vssd1 vccd1 vccd1 _08566_ sky130_fd_sc_hd__or2b_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14903_ _07512_ _07516_ vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__nor2_4
XTAP_5363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18671_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.wall_tracer.rayAddendY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__or2_1
X_15883_ _08493_ _08494_ _08495_ vssd1 vssd1 vccd1 vccd1 _08497_ sky130_fd_sc_hd__a21o_1
XTAP_5385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17622_ _10087_ _10153_ _10157_ vssd1 vssd1 vccd1 vccd1 _10158_ sky130_fd_sc_hd__a21oi_1
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14834_ _07099_ _07195_ _07198_ vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__and3_1
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17553_ _10048_ _10089_ vssd1 vssd1 vccd1 vccd1 _10090_ sky130_fd_sc_hd__xnor2_1
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14765_ _07378_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__clkbuf_4
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11977_ _04665_ o_rgb[14] vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__or2_1
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16504_ _08629_ _04938_ rbzero.wall_tracer.visualWallDist\[11\] vssd1 vssd1 vccd1
+ vccd1 _09113_ sky130_fd_sc_hd__or3b_1
XFILLER_186_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13716_ _06385_ _06393_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__xnor2_2
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17484_ _09762_ _10021_ vssd1 vssd1 vccd1 vccd1 _10022_ sky130_fd_sc_hd__nand2_1
XFILLER_205_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10928_ rbzero.tex_b0\[34\] rbzero.tex_b0\[33\] _03682_ vssd1 vssd1 vccd1 vccd1 _03691_
+ sky130_fd_sc_hd__mux2_1
X_14696_ _07322_ vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19223_ _02786_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__inv_2
X_16435_ _09043_ _09044_ vssd1 vssd1 vccd1 vccd1 _09045_ sky130_fd_sc_hd__nand2_1
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13647_ _06308_ _06322_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__nand2_1
XFILLER_220_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10859_ rbzero.tex_g0\[3\] rbzero.tex_g0\[2\] _03649_ vssd1 vssd1 vccd1 vccd1 _03655_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19154_ rbzero.floor_leak\[4\] _02744_ _02750_ _02738_ vssd1 vssd1 vccd1 vccd1 _00747_
+ sky130_fd_sc_hd__o211a_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _08885_ _08901_ vssd1 vssd1 vccd1 vccd1 _08976_ sky130_fd_sc_hd__nand2_1
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _05434_ _06266_ _05848_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__or3_1
XFILLER_201_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18105_ _01871_ _01885_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15317_ _07783_ _07812_ vssd1 vssd1 vccd1 vccd1 _07931_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12529_ _03789_ _05215_ _05216_ _05217_ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__o2bb2a_2
X_19085_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[2\] _02703_
+ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__mux2_1
X_16297_ _07858_ _07817_ vssd1 vssd1 vccd1 vccd1 _08908_ sky130_fd_sc_hd__nor2_1
XFILLER_157_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18036_ _01728_ _01729_ _01817_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__a21oi_1
XFILLER_117_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15248_ _07400_ _07712_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__nor2_1
XFILLER_133_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15179_ _07519_ _07491_ _07495_ _07500_ vssd1 vssd1 vccd1 vccd1 _07793_ sky130_fd_sc_hd__a31o_2
XFILLER_154_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19987_ _03121_ vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__clkinv_2
XFILLER_101_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18938_ rbzero.pov.spi_buffer\[18\] rbzero.pov.ready_buffer\[18\] _02618_ vssd1 vssd1
+ vccd1 vccd1 _02628_ sky130_fd_sc_hd__mux2_1
.ends

