// This is the unpowered netlist.
module top_ew_algofoogle (i_clk,
    i_debug_map_overlay,
    i_debug_trace_overlay,
    i_debug_vec_overlay,
    i_reg_csb,
    i_reg_mosi,
    i_reg_sclk,
    i_reset_lock_a,
    i_reset_lock_b,
    i_vec_csb,
    i_vec_mosi,
    i_vec_sclk,
    o_hsync,
    o_tex_csb,
    o_tex_oeb0,
    o_tex_out0,
    o_tex_sclk,
    o_vsync,
    i_gpout0_sel,
    i_gpout1_sel,
    i_gpout2_sel,
    i_gpout3_sel,
    i_gpout4_sel,
    i_gpout5_sel,
    i_mode,
    i_tex_in,
    o_gpout,
    o_rgb);
 input i_clk;
 input i_debug_map_overlay;
 input i_debug_trace_overlay;
 input i_debug_vec_overlay;
 input i_reg_csb;
 input i_reg_mosi;
 input i_reg_sclk;
 input i_reset_lock_a;
 input i_reset_lock_b;
 input i_vec_csb;
 input i_vec_mosi;
 input i_vec_sclk;
 output o_hsync;
 output o_tex_csb;
 output o_tex_oeb0;
 output o_tex_out0;
 output o_tex_sclk;
 output o_vsync;
 input [5:0] i_gpout0_sel;
 input [5:0] i_gpout1_sel;
 input [5:0] i_gpout2_sel;
 input [5:0] i_gpout3_sel;
 input [5:0] i_gpout4_sel;
 input [5:0] i_gpout5_sel;
 input [2:0] i_mode;
 input [3:0] i_tex_in;
 output [5:0] o_gpout;
 output [23:0] o_rgb;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire \gpout0.clk_div[0] ;
 wire \gpout0.clk_div[1] ;
 wire \gpout0.hpos[0] ;
 wire \gpout0.hpos[1] ;
 wire \gpout0.hpos[2] ;
 wire \gpout0.hpos[3] ;
 wire \gpout0.hpos[4] ;
 wire \gpout0.hpos[5] ;
 wire \gpout0.hpos[6] ;
 wire \gpout0.hpos[7] ;
 wire \gpout0.hpos[8] ;
 wire \gpout0.hpos[9] ;
 wire \gpout0.vpos[0] ;
 wire \gpout0.vpos[1] ;
 wire \gpout0.vpos[2] ;
 wire \gpout0.vpos[3] ;
 wire \gpout0.vpos[4] ;
 wire \gpout0.vpos[5] ;
 wire \gpout0.vpos[6] ;
 wire \gpout0.vpos[7] ;
 wire \gpout0.vpos[8] ;
 wire \gpout0.vpos[9] ;
 wire \gpout1.clk_div[0] ;
 wire \gpout1.clk_div[1] ;
 wire \gpout2.clk_div[0] ;
 wire \gpout2.clk_div[1] ;
 wire \gpout3.clk_div[0] ;
 wire \gpout3.clk_div[1] ;
 wire \gpout4.clk_div[0] ;
 wire \gpout4.clk_div[1] ;
 wire \gpout5.clk_div[0] ;
 wire \gpout5.clk_div[1] ;
 wire net143;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net144;
 wire net159;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire \rbzero.color_floor[0] ;
 wire \rbzero.color_floor[1] ;
 wire \rbzero.color_floor[2] ;
 wire \rbzero.color_floor[3] ;
 wire \rbzero.color_floor[4] ;
 wire \rbzero.color_floor[5] ;
 wire \rbzero.color_sky[0] ;
 wire \rbzero.color_sky[1] ;
 wire \rbzero.color_sky[2] ;
 wire \rbzero.color_sky[3] ;
 wire \rbzero.color_sky[4] ;
 wire \rbzero.color_sky[5] ;
 wire \rbzero.debug_overlay.facingX[-1] ;
 wire \rbzero.debug_overlay.facingX[-2] ;
 wire \rbzero.debug_overlay.facingX[-3] ;
 wire \rbzero.debug_overlay.facingX[-4] ;
 wire \rbzero.debug_overlay.facingX[-5] ;
 wire \rbzero.debug_overlay.facingX[-6] ;
 wire \rbzero.debug_overlay.facingX[-7] ;
 wire \rbzero.debug_overlay.facingX[-8] ;
 wire \rbzero.debug_overlay.facingX[-9] ;
 wire \rbzero.debug_overlay.facingX[0] ;
 wire \rbzero.debug_overlay.facingX[10] ;
 wire \rbzero.debug_overlay.facingY[-1] ;
 wire \rbzero.debug_overlay.facingY[-2] ;
 wire \rbzero.debug_overlay.facingY[-3] ;
 wire \rbzero.debug_overlay.facingY[-4] ;
 wire \rbzero.debug_overlay.facingY[-5] ;
 wire \rbzero.debug_overlay.facingY[-6] ;
 wire \rbzero.debug_overlay.facingY[-7] ;
 wire \rbzero.debug_overlay.facingY[-8] ;
 wire \rbzero.debug_overlay.facingY[-9] ;
 wire \rbzero.debug_overlay.facingY[0] ;
 wire \rbzero.debug_overlay.facingY[10] ;
 wire \rbzero.debug_overlay.playerX[-1] ;
 wire \rbzero.debug_overlay.playerX[-2] ;
 wire \rbzero.debug_overlay.playerX[-3] ;
 wire \rbzero.debug_overlay.playerX[-4] ;
 wire \rbzero.debug_overlay.playerX[-5] ;
 wire \rbzero.debug_overlay.playerX[-6] ;
 wire \rbzero.debug_overlay.playerX[-7] ;
 wire \rbzero.debug_overlay.playerX[-8] ;
 wire \rbzero.debug_overlay.playerX[-9] ;
 wire \rbzero.debug_overlay.playerX[0] ;
 wire \rbzero.debug_overlay.playerX[1] ;
 wire \rbzero.debug_overlay.playerX[2] ;
 wire \rbzero.debug_overlay.playerX[3] ;
 wire \rbzero.debug_overlay.playerX[4] ;
 wire \rbzero.debug_overlay.playerX[5] ;
 wire \rbzero.debug_overlay.playerY[-1] ;
 wire \rbzero.debug_overlay.playerY[-2] ;
 wire \rbzero.debug_overlay.playerY[-3] ;
 wire \rbzero.debug_overlay.playerY[-4] ;
 wire \rbzero.debug_overlay.playerY[-5] ;
 wire \rbzero.debug_overlay.playerY[-6] ;
 wire \rbzero.debug_overlay.playerY[-7] ;
 wire \rbzero.debug_overlay.playerY[-8] ;
 wire \rbzero.debug_overlay.playerY[-9] ;
 wire \rbzero.debug_overlay.playerY[0] ;
 wire \rbzero.debug_overlay.playerY[1] ;
 wire \rbzero.debug_overlay.playerY[2] ;
 wire \rbzero.debug_overlay.playerY[3] ;
 wire \rbzero.debug_overlay.playerY[4] ;
 wire \rbzero.debug_overlay.playerY[5] ;
 wire \rbzero.debug_overlay.vplaneX[-1] ;
 wire \rbzero.debug_overlay.vplaneX[-2] ;
 wire \rbzero.debug_overlay.vplaneX[-3] ;
 wire \rbzero.debug_overlay.vplaneX[-4] ;
 wire \rbzero.debug_overlay.vplaneX[-5] ;
 wire \rbzero.debug_overlay.vplaneX[-6] ;
 wire \rbzero.debug_overlay.vplaneX[-7] ;
 wire \rbzero.debug_overlay.vplaneX[-8] ;
 wire \rbzero.debug_overlay.vplaneX[-9] ;
 wire \rbzero.debug_overlay.vplaneX[0] ;
 wire \rbzero.debug_overlay.vplaneX[10] ;
 wire \rbzero.debug_overlay.vplaneY[-1] ;
 wire \rbzero.debug_overlay.vplaneY[-2] ;
 wire \rbzero.debug_overlay.vplaneY[-3] ;
 wire \rbzero.debug_overlay.vplaneY[-4] ;
 wire \rbzero.debug_overlay.vplaneY[-5] ;
 wire \rbzero.debug_overlay.vplaneY[-6] ;
 wire \rbzero.debug_overlay.vplaneY[-7] ;
 wire \rbzero.debug_overlay.vplaneY[-8] ;
 wire \rbzero.debug_overlay.vplaneY[-9] ;
 wire \rbzero.debug_overlay.vplaneY[0] ;
 wire \rbzero.debug_overlay.vplaneY[10] ;
 wire \rbzero.floor_leak[0] ;
 wire \rbzero.floor_leak[1] ;
 wire \rbzero.floor_leak[2] ;
 wire \rbzero.floor_leak[3] ;
 wire \rbzero.floor_leak[4] ;
 wire \rbzero.floor_leak[5] ;
 wire \rbzero.hsync ;
 wire \rbzero.map_rom.a6 ;
 wire \rbzero.map_rom.b6 ;
 wire \rbzero.map_rom.c6 ;
 wire \rbzero.map_rom.d6 ;
 wire \rbzero.map_rom.f1 ;
 wire \rbzero.map_rom.f2 ;
 wire \rbzero.map_rom.f3 ;
 wire \rbzero.map_rom.f4 ;
 wire \rbzero.map_rom.i_col[4] ;
 wire \rbzero.map_rom.i_row[4] ;
 wire \rbzero.otherx[0] ;
 wire \rbzero.otherx[1] ;
 wire \rbzero.otherx[2] ;
 wire \rbzero.otherx[3] ;
 wire \rbzero.otherx[4] ;
 wire \rbzero.othery[0] ;
 wire \rbzero.othery[1] ;
 wire \rbzero.othery[2] ;
 wire \rbzero.othery[3] ;
 wire \rbzero.othery[4] ;
 wire \rbzero.pov.mosi ;
 wire \rbzero.pov.mosi_buffer[0] ;
 wire \rbzero.pov.ready ;
 wire \rbzero.pov.ready_buffer[0] ;
 wire \rbzero.pov.ready_buffer[10] ;
 wire \rbzero.pov.ready_buffer[11] ;
 wire \rbzero.pov.ready_buffer[12] ;
 wire \rbzero.pov.ready_buffer[13] ;
 wire \rbzero.pov.ready_buffer[14] ;
 wire \rbzero.pov.ready_buffer[15] ;
 wire \rbzero.pov.ready_buffer[16] ;
 wire \rbzero.pov.ready_buffer[17] ;
 wire \rbzero.pov.ready_buffer[18] ;
 wire \rbzero.pov.ready_buffer[19] ;
 wire \rbzero.pov.ready_buffer[1] ;
 wire \rbzero.pov.ready_buffer[20] ;
 wire \rbzero.pov.ready_buffer[21] ;
 wire \rbzero.pov.ready_buffer[22] ;
 wire \rbzero.pov.ready_buffer[23] ;
 wire \rbzero.pov.ready_buffer[24] ;
 wire \rbzero.pov.ready_buffer[25] ;
 wire \rbzero.pov.ready_buffer[26] ;
 wire \rbzero.pov.ready_buffer[27] ;
 wire \rbzero.pov.ready_buffer[28] ;
 wire \rbzero.pov.ready_buffer[29] ;
 wire \rbzero.pov.ready_buffer[2] ;
 wire \rbzero.pov.ready_buffer[30] ;
 wire \rbzero.pov.ready_buffer[31] ;
 wire \rbzero.pov.ready_buffer[32] ;
 wire \rbzero.pov.ready_buffer[33] ;
 wire \rbzero.pov.ready_buffer[34] ;
 wire \rbzero.pov.ready_buffer[35] ;
 wire \rbzero.pov.ready_buffer[36] ;
 wire \rbzero.pov.ready_buffer[37] ;
 wire \rbzero.pov.ready_buffer[38] ;
 wire \rbzero.pov.ready_buffer[39] ;
 wire \rbzero.pov.ready_buffer[3] ;
 wire \rbzero.pov.ready_buffer[40] ;
 wire \rbzero.pov.ready_buffer[41] ;
 wire \rbzero.pov.ready_buffer[42] ;
 wire \rbzero.pov.ready_buffer[43] ;
 wire \rbzero.pov.ready_buffer[44] ;
 wire \rbzero.pov.ready_buffer[45] ;
 wire \rbzero.pov.ready_buffer[46] ;
 wire \rbzero.pov.ready_buffer[47] ;
 wire \rbzero.pov.ready_buffer[48] ;
 wire \rbzero.pov.ready_buffer[49] ;
 wire \rbzero.pov.ready_buffer[4] ;
 wire \rbzero.pov.ready_buffer[50] ;
 wire \rbzero.pov.ready_buffer[51] ;
 wire \rbzero.pov.ready_buffer[52] ;
 wire \rbzero.pov.ready_buffer[53] ;
 wire \rbzero.pov.ready_buffer[54] ;
 wire \rbzero.pov.ready_buffer[55] ;
 wire \rbzero.pov.ready_buffer[56] ;
 wire \rbzero.pov.ready_buffer[57] ;
 wire \rbzero.pov.ready_buffer[58] ;
 wire \rbzero.pov.ready_buffer[59] ;
 wire \rbzero.pov.ready_buffer[5] ;
 wire \rbzero.pov.ready_buffer[60] ;
 wire \rbzero.pov.ready_buffer[61] ;
 wire \rbzero.pov.ready_buffer[62] ;
 wire \rbzero.pov.ready_buffer[63] ;
 wire \rbzero.pov.ready_buffer[64] ;
 wire \rbzero.pov.ready_buffer[65] ;
 wire \rbzero.pov.ready_buffer[66] ;
 wire \rbzero.pov.ready_buffer[67] ;
 wire \rbzero.pov.ready_buffer[68] ;
 wire \rbzero.pov.ready_buffer[69] ;
 wire \rbzero.pov.ready_buffer[6] ;
 wire \rbzero.pov.ready_buffer[70] ;
 wire \rbzero.pov.ready_buffer[71] ;
 wire \rbzero.pov.ready_buffer[72] ;
 wire \rbzero.pov.ready_buffer[73] ;
 wire \rbzero.pov.ready_buffer[7] ;
 wire \rbzero.pov.ready_buffer[8] ;
 wire \rbzero.pov.ready_buffer[9] ;
 wire \rbzero.pov.sclk_buffer[0] ;
 wire \rbzero.pov.sclk_buffer[1] ;
 wire \rbzero.pov.sclk_buffer[2] ;
 wire \rbzero.pov.spi_buffer[0] ;
 wire \rbzero.pov.spi_buffer[10] ;
 wire \rbzero.pov.spi_buffer[11] ;
 wire \rbzero.pov.spi_buffer[12] ;
 wire \rbzero.pov.spi_buffer[13] ;
 wire \rbzero.pov.spi_buffer[14] ;
 wire \rbzero.pov.spi_buffer[15] ;
 wire \rbzero.pov.spi_buffer[16] ;
 wire \rbzero.pov.spi_buffer[17] ;
 wire \rbzero.pov.spi_buffer[18] ;
 wire \rbzero.pov.spi_buffer[19] ;
 wire \rbzero.pov.spi_buffer[1] ;
 wire \rbzero.pov.spi_buffer[20] ;
 wire \rbzero.pov.spi_buffer[21] ;
 wire \rbzero.pov.spi_buffer[22] ;
 wire \rbzero.pov.spi_buffer[23] ;
 wire \rbzero.pov.spi_buffer[24] ;
 wire \rbzero.pov.spi_buffer[25] ;
 wire \rbzero.pov.spi_buffer[26] ;
 wire \rbzero.pov.spi_buffer[27] ;
 wire \rbzero.pov.spi_buffer[28] ;
 wire \rbzero.pov.spi_buffer[29] ;
 wire \rbzero.pov.spi_buffer[2] ;
 wire \rbzero.pov.spi_buffer[30] ;
 wire \rbzero.pov.spi_buffer[31] ;
 wire \rbzero.pov.spi_buffer[32] ;
 wire \rbzero.pov.spi_buffer[33] ;
 wire \rbzero.pov.spi_buffer[34] ;
 wire \rbzero.pov.spi_buffer[35] ;
 wire \rbzero.pov.spi_buffer[36] ;
 wire \rbzero.pov.spi_buffer[37] ;
 wire \rbzero.pov.spi_buffer[38] ;
 wire \rbzero.pov.spi_buffer[39] ;
 wire \rbzero.pov.spi_buffer[3] ;
 wire \rbzero.pov.spi_buffer[40] ;
 wire \rbzero.pov.spi_buffer[41] ;
 wire \rbzero.pov.spi_buffer[42] ;
 wire \rbzero.pov.spi_buffer[43] ;
 wire \rbzero.pov.spi_buffer[44] ;
 wire \rbzero.pov.spi_buffer[45] ;
 wire \rbzero.pov.spi_buffer[46] ;
 wire \rbzero.pov.spi_buffer[47] ;
 wire \rbzero.pov.spi_buffer[48] ;
 wire \rbzero.pov.spi_buffer[49] ;
 wire \rbzero.pov.spi_buffer[4] ;
 wire \rbzero.pov.spi_buffer[50] ;
 wire \rbzero.pov.spi_buffer[51] ;
 wire \rbzero.pov.spi_buffer[52] ;
 wire \rbzero.pov.spi_buffer[53] ;
 wire \rbzero.pov.spi_buffer[54] ;
 wire \rbzero.pov.spi_buffer[55] ;
 wire \rbzero.pov.spi_buffer[56] ;
 wire \rbzero.pov.spi_buffer[57] ;
 wire \rbzero.pov.spi_buffer[58] ;
 wire \rbzero.pov.spi_buffer[59] ;
 wire \rbzero.pov.spi_buffer[5] ;
 wire \rbzero.pov.spi_buffer[60] ;
 wire \rbzero.pov.spi_buffer[61] ;
 wire \rbzero.pov.spi_buffer[62] ;
 wire \rbzero.pov.spi_buffer[63] ;
 wire \rbzero.pov.spi_buffer[64] ;
 wire \rbzero.pov.spi_buffer[65] ;
 wire \rbzero.pov.spi_buffer[66] ;
 wire \rbzero.pov.spi_buffer[67] ;
 wire \rbzero.pov.spi_buffer[68] ;
 wire \rbzero.pov.spi_buffer[69] ;
 wire \rbzero.pov.spi_buffer[6] ;
 wire \rbzero.pov.spi_buffer[70] ;
 wire \rbzero.pov.spi_buffer[71] ;
 wire \rbzero.pov.spi_buffer[72] ;
 wire \rbzero.pov.spi_buffer[73] ;
 wire \rbzero.pov.spi_buffer[7] ;
 wire \rbzero.pov.spi_buffer[8] ;
 wire \rbzero.pov.spi_buffer[9] ;
 wire \rbzero.pov.spi_counter[0] ;
 wire \rbzero.pov.spi_counter[1] ;
 wire \rbzero.pov.spi_counter[2] ;
 wire \rbzero.pov.spi_counter[3] ;
 wire \rbzero.pov.spi_counter[4] ;
 wire \rbzero.pov.spi_counter[5] ;
 wire \rbzero.pov.spi_counter[6] ;
 wire \rbzero.pov.spi_done ;
 wire \rbzero.pov.ss_buffer[0] ;
 wire \rbzero.pov.ss_buffer[1] ;
 wire \rbzero.row_render.side ;
 wire \rbzero.row_render.size[0] ;
 wire \rbzero.row_render.size[10] ;
 wire \rbzero.row_render.size[1] ;
 wire \rbzero.row_render.size[2] ;
 wire \rbzero.row_render.size[3] ;
 wire \rbzero.row_render.size[4] ;
 wire \rbzero.row_render.size[5] ;
 wire \rbzero.row_render.size[6] ;
 wire \rbzero.row_render.size[7] ;
 wire \rbzero.row_render.size[8] ;
 wire \rbzero.row_render.size[9] ;
 wire \rbzero.row_render.texu[0] ;
 wire \rbzero.row_render.texu[1] ;
 wire \rbzero.row_render.texu[2] ;
 wire \rbzero.row_render.texu[3] ;
 wire \rbzero.row_render.texu[4] ;
 wire \rbzero.row_render.texu[5] ;
 wire \rbzero.row_render.vinf ;
 wire \rbzero.row_render.wall[0] ;
 wire \rbzero.row_render.wall[1] ;
 wire \rbzero.spi_registers.got_new_floor ;
 wire \rbzero.spi_registers.got_new_leak ;
 wire \rbzero.spi_registers.got_new_other ;
 wire \rbzero.spi_registers.got_new_sky ;
 wire \rbzero.spi_registers.got_new_vinf ;
 wire \rbzero.spi_registers.got_new_vshift ;
 wire \rbzero.spi_registers.mosi ;
 wire \rbzero.spi_registers.mosi_buffer[0] ;
 wire \rbzero.spi_registers.new_floor[0] ;
 wire \rbzero.spi_registers.new_floor[1] ;
 wire \rbzero.spi_registers.new_floor[2] ;
 wire \rbzero.spi_registers.new_floor[3] ;
 wire \rbzero.spi_registers.new_floor[4] ;
 wire \rbzero.spi_registers.new_floor[5] ;
 wire \rbzero.spi_registers.new_leak[0] ;
 wire \rbzero.spi_registers.new_leak[1] ;
 wire \rbzero.spi_registers.new_leak[2] ;
 wire \rbzero.spi_registers.new_leak[3] ;
 wire \rbzero.spi_registers.new_leak[4] ;
 wire \rbzero.spi_registers.new_leak[5] ;
 wire \rbzero.spi_registers.new_other[0] ;
 wire \rbzero.spi_registers.new_other[10] ;
 wire \rbzero.spi_registers.new_other[1] ;
 wire \rbzero.spi_registers.new_other[2] ;
 wire \rbzero.spi_registers.new_other[3] ;
 wire \rbzero.spi_registers.new_other[4] ;
 wire \rbzero.spi_registers.new_other[6] ;
 wire \rbzero.spi_registers.new_other[7] ;
 wire \rbzero.spi_registers.new_other[8] ;
 wire \rbzero.spi_registers.new_other[9] ;
 wire \rbzero.spi_registers.new_sky[0] ;
 wire \rbzero.spi_registers.new_sky[1] ;
 wire \rbzero.spi_registers.new_sky[2] ;
 wire \rbzero.spi_registers.new_sky[3] ;
 wire \rbzero.spi_registers.new_sky[4] ;
 wire \rbzero.spi_registers.new_sky[5] ;
 wire \rbzero.spi_registers.new_vinf ;
 wire \rbzero.spi_registers.new_vshift[0] ;
 wire \rbzero.spi_registers.new_vshift[1] ;
 wire \rbzero.spi_registers.new_vshift[2] ;
 wire \rbzero.spi_registers.new_vshift[3] ;
 wire \rbzero.spi_registers.new_vshift[4] ;
 wire \rbzero.spi_registers.new_vshift[5] ;
 wire \rbzero.spi_registers.sclk_buffer[0] ;
 wire \rbzero.spi_registers.sclk_buffer[1] ;
 wire \rbzero.spi_registers.sclk_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[0] ;
 wire \rbzero.spi_registers.spi_buffer[10] ;
 wire \rbzero.spi_registers.spi_buffer[1] ;
 wire \rbzero.spi_registers.spi_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[3] ;
 wire \rbzero.spi_registers.spi_buffer[4] ;
 wire \rbzero.spi_registers.spi_buffer[5] ;
 wire \rbzero.spi_registers.spi_buffer[6] ;
 wire \rbzero.spi_registers.spi_buffer[7] ;
 wire \rbzero.spi_registers.spi_buffer[8] ;
 wire \rbzero.spi_registers.spi_buffer[9] ;
 wire \rbzero.spi_registers.spi_cmd[0] ;
 wire \rbzero.spi_registers.spi_cmd[1] ;
 wire \rbzero.spi_registers.spi_cmd[2] ;
 wire \rbzero.spi_registers.spi_cmd[3] ;
 wire \rbzero.spi_registers.spi_counter[0] ;
 wire \rbzero.spi_registers.spi_counter[1] ;
 wire \rbzero.spi_registers.spi_counter[2] ;
 wire \rbzero.spi_registers.spi_counter[3] ;
 wire \rbzero.spi_registers.spi_counter[4] ;
 wire \rbzero.spi_registers.spi_counter[5] ;
 wire \rbzero.spi_registers.spi_counter[6] ;
 wire \rbzero.spi_registers.spi_done ;
 wire \rbzero.spi_registers.ss_buffer[0] ;
 wire \rbzero.spi_registers.ss_buffer[1] ;
 wire \rbzero.spi_registers.vshift[0] ;
 wire \rbzero.spi_registers.vshift[1] ;
 wire \rbzero.spi_registers.vshift[2] ;
 wire \rbzero.spi_registers.vshift[3] ;
 wire \rbzero.spi_registers.vshift[4] ;
 wire \rbzero.spi_registers.vshift[5] ;
 wire \rbzero.texV[-10] ;
 wire \rbzero.texV[-11] ;
 wire \rbzero.texV[-12] ;
 wire \rbzero.texV[-1] ;
 wire \rbzero.texV[-2] ;
 wire \rbzero.texV[-3] ;
 wire \rbzero.texV[-4] ;
 wire \rbzero.texV[-5] ;
 wire \rbzero.texV[-6] ;
 wire \rbzero.texV[-7] ;
 wire \rbzero.texV[-8] ;
 wire \rbzero.texV[-9] ;
 wire \rbzero.texV[0] ;
 wire \rbzero.texV[10] ;
 wire \rbzero.texV[11] ;
 wire \rbzero.texV[1] ;
 wire \rbzero.texV[2] ;
 wire \rbzero.texV[3] ;
 wire \rbzero.texV[4] ;
 wire \rbzero.texV[5] ;
 wire \rbzero.texV[6] ;
 wire \rbzero.texV[7] ;
 wire \rbzero.texV[8] ;
 wire \rbzero.texV[9] ;
 wire \rbzero.tex_b0[0] ;
 wire \rbzero.tex_b0[10] ;
 wire \rbzero.tex_b0[11] ;
 wire \rbzero.tex_b0[12] ;
 wire \rbzero.tex_b0[13] ;
 wire \rbzero.tex_b0[14] ;
 wire \rbzero.tex_b0[15] ;
 wire \rbzero.tex_b0[16] ;
 wire \rbzero.tex_b0[17] ;
 wire \rbzero.tex_b0[18] ;
 wire \rbzero.tex_b0[19] ;
 wire \rbzero.tex_b0[1] ;
 wire \rbzero.tex_b0[20] ;
 wire \rbzero.tex_b0[21] ;
 wire \rbzero.tex_b0[22] ;
 wire \rbzero.tex_b0[23] ;
 wire \rbzero.tex_b0[24] ;
 wire \rbzero.tex_b0[25] ;
 wire \rbzero.tex_b0[26] ;
 wire \rbzero.tex_b0[27] ;
 wire \rbzero.tex_b0[28] ;
 wire \rbzero.tex_b0[29] ;
 wire \rbzero.tex_b0[2] ;
 wire \rbzero.tex_b0[30] ;
 wire \rbzero.tex_b0[31] ;
 wire \rbzero.tex_b0[32] ;
 wire \rbzero.tex_b0[33] ;
 wire \rbzero.tex_b0[34] ;
 wire \rbzero.tex_b0[35] ;
 wire \rbzero.tex_b0[36] ;
 wire \rbzero.tex_b0[37] ;
 wire \rbzero.tex_b0[38] ;
 wire \rbzero.tex_b0[39] ;
 wire \rbzero.tex_b0[3] ;
 wire \rbzero.tex_b0[40] ;
 wire \rbzero.tex_b0[41] ;
 wire \rbzero.tex_b0[42] ;
 wire \rbzero.tex_b0[43] ;
 wire \rbzero.tex_b0[44] ;
 wire \rbzero.tex_b0[45] ;
 wire \rbzero.tex_b0[46] ;
 wire \rbzero.tex_b0[47] ;
 wire \rbzero.tex_b0[48] ;
 wire \rbzero.tex_b0[49] ;
 wire \rbzero.tex_b0[4] ;
 wire \rbzero.tex_b0[50] ;
 wire \rbzero.tex_b0[51] ;
 wire \rbzero.tex_b0[52] ;
 wire \rbzero.tex_b0[53] ;
 wire \rbzero.tex_b0[54] ;
 wire \rbzero.tex_b0[55] ;
 wire \rbzero.tex_b0[56] ;
 wire \rbzero.tex_b0[57] ;
 wire \rbzero.tex_b0[58] ;
 wire \rbzero.tex_b0[59] ;
 wire \rbzero.tex_b0[5] ;
 wire \rbzero.tex_b0[60] ;
 wire \rbzero.tex_b0[61] ;
 wire \rbzero.tex_b0[62] ;
 wire \rbzero.tex_b0[63] ;
 wire \rbzero.tex_b0[6] ;
 wire \rbzero.tex_b0[7] ;
 wire \rbzero.tex_b0[8] ;
 wire \rbzero.tex_b0[9] ;
 wire \rbzero.tex_b1[0] ;
 wire \rbzero.tex_b1[10] ;
 wire \rbzero.tex_b1[11] ;
 wire \rbzero.tex_b1[12] ;
 wire \rbzero.tex_b1[13] ;
 wire \rbzero.tex_b1[14] ;
 wire \rbzero.tex_b1[15] ;
 wire \rbzero.tex_b1[16] ;
 wire \rbzero.tex_b1[17] ;
 wire \rbzero.tex_b1[18] ;
 wire \rbzero.tex_b1[19] ;
 wire \rbzero.tex_b1[1] ;
 wire \rbzero.tex_b1[20] ;
 wire \rbzero.tex_b1[21] ;
 wire \rbzero.tex_b1[22] ;
 wire \rbzero.tex_b1[23] ;
 wire \rbzero.tex_b1[24] ;
 wire \rbzero.tex_b1[25] ;
 wire \rbzero.tex_b1[26] ;
 wire \rbzero.tex_b1[27] ;
 wire \rbzero.tex_b1[28] ;
 wire \rbzero.tex_b1[29] ;
 wire \rbzero.tex_b1[2] ;
 wire \rbzero.tex_b1[30] ;
 wire \rbzero.tex_b1[31] ;
 wire \rbzero.tex_b1[32] ;
 wire \rbzero.tex_b1[33] ;
 wire \rbzero.tex_b1[34] ;
 wire \rbzero.tex_b1[35] ;
 wire \rbzero.tex_b1[36] ;
 wire \rbzero.tex_b1[37] ;
 wire \rbzero.tex_b1[38] ;
 wire \rbzero.tex_b1[39] ;
 wire \rbzero.tex_b1[3] ;
 wire \rbzero.tex_b1[40] ;
 wire \rbzero.tex_b1[41] ;
 wire \rbzero.tex_b1[42] ;
 wire \rbzero.tex_b1[43] ;
 wire \rbzero.tex_b1[44] ;
 wire \rbzero.tex_b1[45] ;
 wire \rbzero.tex_b1[46] ;
 wire \rbzero.tex_b1[47] ;
 wire \rbzero.tex_b1[48] ;
 wire \rbzero.tex_b1[49] ;
 wire \rbzero.tex_b1[4] ;
 wire \rbzero.tex_b1[50] ;
 wire \rbzero.tex_b1[51] ;
 wire \rbzero.tex_b1[52] ;
 wire \rbzero.tex_b1[53] ;
 wire \rbzero.tex_b1[54] ;
 wire \rbzero.tex_b1[55] ;
 wire \rbzero.tex_b1[56] ;
 wire \rbzero.tex_b1[57] ;
 wire \rbzero.tex_b1[58] ;
 wire \rbzero.tex_b1[59] ;
 wire \rbzero.tex_b1[5] ;
 wire \rbzero.tex_b1[60] ;
 wire \rbzero.tex_b1[61] ;
 wire \rbzero.tex_b1[62] ;
 wire \rbzero.tex_b1[63] ;
 wire \rbzero.tex_b1[6] ;
 wire \rbzero.tex_b1[7] ;
 wire \rbzero.tex_b1[8] ;
 wire \rbzero.tex_b1[9] ;
 wire \rbzero.tex_g0[0] ;
 wire \rbzero.tex_g0[10] ;
 wire \rbzero.tex_g0[11] ;
 wire \rbzero.tex_g0[12] ;
 wire \rbzero.tex_g0[13] ;
 wire \rbzero.tex_g0[14] ;
 wire \rbzero.tex_g0[15] ;
 wire \rbzero.tex_g0[16] ;
 wire \rbzero.tex_g0[17] ;
 wire \rbzero.tex_g0[18] ;
 wire \rbzero.tex_g0[19] ;
 wire \rbzero.tex_g0[1] ;
 wire \rbzero.tex_g0[20] ;
 wire \rbzero.tex_g0[21] ;
 wire \rbzero.tex_g0[22] ;
 wire \rbzero.tex_g0[23] ;
 wire \rbzero.tex_g0[24] ;
 wire \rbzero.tex_g0[25] ;
 wire \rbzero.tex_g0[26] ;
 wire \rbzero.tex_g0[27] ;
 wire \rbzero.tex_g0[28] ;
 wire \rbzero.tex_g0[29] ;
 wire \rbzero.tex_g0[2] ;
 wire \rbzero.tex_g0[30] ;
 wire \rbzero.tex_g0[31] ;
 wire \rbzero.tex_g0[32] ;
 wire \rbzero.tex_g0[33] ;
 wire \rbzero.tex_g0[34] ;
 wire \rbzero.tex_g0[35] ;
 wire \rbzero.tex_g0[36] ;
 wire \rbzero.tex_g0[37] ;
 wire \rbzero.tex_g0[38] ;
 wire \rbzero.tex_g0[39] ;
 wire \rbzero.tex_g0[3] ;
 wire \rbzero.tex_g0[40] ;
 wire \rbzero.tex_g0[41] ;
 wire \rbzero.tex_g0[42] ;
 wire \rbzero.tex_g0[43] ;
 wire \rbzero.tex_g0[44] ;
 wire \rbzero.tex_g0[45] ;
 wire \rbzero.tex_g0[46] ;
 wire \rbzero.tex_g0[47] ;
 wire \rbzero.tex_g0[48] ;
 wire \rbzero.tex_g0[49] ;
 wire \rbzero.tex_g0[4] ;
 wire \rbzero.tex_g0[50] ;
 wire \rbzero.tex_g0[51] ;
 wire \rbzero.tex_g0[52] ;
 wire \rbzero.tex_g0[53] ;
 wire \rbzero.tex_g0[54] ;
 wire \rbzero.tex_g0[55] ;
 wire \rbzero.tex_g0[56] ;
 wire \rbzero.tex_g0[57] ;
 wire \rbzero.tex_g0[58] ;
 wire \rbzero.tex_g0[59] ;
 wire \rbzero.tex_g0[5] ;
 wire \rbzero.tex_g0[60] ;
 wire \rbzero.tex_g0[61] ;
 wire \rbzero.tex_g0[62] ;
 wire \rbzero.tex_g0[63] ;
 wire \rbzero.tex_g0[6] ;
 wire \rbzero.tex_g0[7] ;
 wire \rbzero.tex_g0[8] ;
 wire \rbzero.tex_g0[9] ;
 wire \rbzero.tex_g1[0] ;
 wire \rbzero.tex_g1[10] ;
 wire \rbzero.tex_g1[11] ;
 wire \rbzero.tex_g1[12] ;
 wire \rbzero.tex_g1[13] ;
 wire \rbzero.tex_g1[14] ;
 wire \rbzero.tex_g1[15] ;
 wire \rbzero.tex_g1[16] ;
 wire \rbzero.tex_g1[17] ;
 wire \rbzero.tex_g1[18] ;
 wire \rbzero.tex_g1[19] ;
 wire \rbzero.tex_g1[1] ;
 wire \rbzero.tex_g1[20] ;
 wire \rbzero.tex_g1[21] ;
 wire \rbzero.tex_g1[22] ;
 wire \rbzero.tex_g1[23] ;
 wire \rbzero.tex_g1[24] ;
 wire \rbzero.tex_g1[25] ;
 wire \rbzero.tex_g1[26] ;
 wire \rbzero.tex_g1[27] ;
 wire \rbzero.tex_g1[28] ;
 wire \rbzero.tex_g1[29] ;
 wire \rbzero.tex_g1[2] ;
 wire \rbzero.tex_g1[30] ;
 wire \rbzero.tex_g1[31] ;
 wire \rbzero.tex_g1[32] ;
 wire \rbzero.tex_g1[33] ;
 wire \rbzero.tex_g1[34] ;
 wire \rbzero.tex_g1[35] ;
 wire \rbzero.tex_g1[36] ;
 wire \rbzero.tex_g1[37] ;
 wire \rbzero.tex_g1[38] ;
 wire \rbzero.tex_g1[39] ;
 wire \rbzero.tex_g1[3] ;
 wire \rbzero.tex_g1[40] ;
 wire \rbzero.tex_g1[41] ;
 wire \rbzero.tex_g1[42] ;
 wire \rbzero.tex_g1[43] ;
 wire \rbzero.tex_g1[44] ;
 wire \rbzero.tex_g1[45] ;
 wire \rbzero.tex_g1[46] ;
 wire \rbzero.tex_g1[47] ;
 wire \rbzero.tex_g1[48] ;
 wire \rbzero.tex_g1[49] ;
 wire \rbzero.tex_g1[4] ;
 wire \rbzero.tex_g1[50] ;
 wire \rbzero.tex_g1[51] ;
 wire \rbzero.tex_g1[52] ;
 wire \rbzero.tex_g1[53] ;
 wire \rbzero.tex_g1[54] ;
 wire \rbzero.tex_g1[55] ;
 wire \rbzero.tex_g1[56] ;
 wire \rbzero.tex_g1[57] ;
 wire \rbzero.tex_g1[58] ;
 wire \rbzero.tex_g1[59] ;
 wire \rbzero.tex_g1[5] ;
 wire \rbzero.tex_g1[60] ;
 wire \rbzero.tex_g1[61] ;
 wire \rbzero.tex_g1[62] ;
 wire \rbzero.tex_g1[63] ;
 wire \rbzero.tex_g1[6] ;
 wire \rbzero.tex_g1[7] ;
 wire \rbzero.tex_g1[8] ;
 wire \rbzero.tex_g1[9] ;
 wire \rbzero.tex_r0[0] ;
 wire \rbzero.tex_r0[10] ;
 wire \rbzero.tex_r0[11] ;
 wire \rbzero.tex_r0[12] ;
 wire \rbzero.tex_r0[13] ;
 wire \rbzero.tex_r0[14] ;
 wire \rbzero.tex_r0[15] ;
 wire \rbzero.tex_r0[16] ;
 wire \rbzero.tex_r0[17] ;
 wire \rbzero.tex_r0[18] ;
 wire \rbzero.tex_r0[19] ;
 wire \rbzero.tex_r0[1] ;
 wire \rbzero.tex_r0[20] ;
 wire \rbzero.tex_r0[21] ;
 wire \rbzero.tex_r0[22] ;
 wire \rbzero.tex_r0[23] ;
 wire \rbzero.tex_r0[24] ;
 wire \rbzero.tex_r0[25] ;
 wire \rbzero.tex_r0[26] ;
 wire \rbzero.tex_r0[27] ;
 wire \rbzero.tex_r0[28] ;
 wire \rbzero.tex_r0[29] ;
 wire \rbzero.tex_r0[2] ;
 wire \rbzero.tex_r0[30] ;
 wire \rbzero.tex_r0[31] ;
 wire \rbzero.tex_r0[32] ;
 wire \rbzero.tex_r0[33] ;
 wire \rbzero.tex_r0[34] ;
 wire \rbzero.tex_r0[35] ;
 wire \rbzero.tex_r0[36] ;
 wire \rbzero.tex_r0[37] ;
 wire \rbzero.tex_r0[38] ;
 wire \rbzero.tex_r0[39] ;
 wire \rbzero.tex_r0[3] ;
 wire \rbzero.tex_r0[40] ;
 wire \rbzero.tex_r0[41] ;
 wire \rbzero.tex_r0[42] ;
 wire \rbzero.tex_r0[43] ;
 wire \rbzero.tex_r0[44] ;
 wire \rbzero.tex_r0[45] ;
 wire \rbzero.tex_r0[46] ;
 wire \rbzero.tex_r0[47] ;
 wire \rbzero.tex_r0[48] ;
 wire \rbzero.tex_r0[49] ;
 wire \rbzero.tex_r0[4] ;
 wire \rbzero.tex_r0[50] ;
 wire \rbzero.tex_r0[51] ;
 wire \rbzero.tex_r0[52] ;
 wire \rbzero.tex_r0[53] ;
 wire \rbzero.tex_r0[54] ;
 wire \rbzero.tex_r0[55] ;
 wire \rbzero.tex_r0[56] ;
 wire \rbzero.tex_r0[57] ;
 wire \rbzero.tex_r0[58] ;
 wire \rbzero.tex_r0[59] ;
 wire \rbzero.tex_r0[5] ;
 wire \rbzero.tex_r0[60] ;
 wire \rbzero.tex_r0[61] ;
 wire \rbzero.tex_r0[62] ;
 wire \rbzero.tex_r0[63] ;
 wire \rbzero.tex_r0[6] ;
 wire \rbzero.tex_r0[7] ;
 wire \rbzero.tex_r0[8] ;
 wire \rbzero.tex_r0[9] ;
 wire \rbzero.tex_r1[0] ;
 wire \rbzero.tex_r1[10] ;
 wire \rbzero.tex_r1[11] ;
 wire \rbzero.tex_r1[12] ;
 wire \rbzero.tex_r1[13] ;
 wire \rbzero.tex_r1[14] ;
 wire \rbzero.tex_r1[15] ;
 wire \rbzero.tex_r1[16] ;
 wire \rbzero.tex_r1[17] ;
 wire \rbzero.tex_r1[18] ;
 wire \rbzero.tex_r1[19] ;
 wire \rbzero.tex_r1[1] ;
 wire \rbzero.tex_r1[20] ;
 wire \rbzero.tex_r1[21] ;
 wire \rbzero.tex_r1[22] ;
 wire \rbzero.tex_r1[23] ;
 wire \rbzero.tex_r1[24] ;
 wire \rbzero.tex_r1[25] ;
 wire \rbzero.tex_r1[26] ;
 wire \rbzero.tex_r1[27] ;
 wire \rbzero.tex_r1[28] ;
 wire \rbzero.tex_r1[29] ;
 wire \rbzero.tex_r1[2] ;
 wire \rbzero.tex_r1[30] ;
 wire \rbzero.tex_r1[31] ;
 wire \rbzero.tex_r1[32] ;
 wire \rbzero.tex_r1[33] ;
 wire \rbzero.tex_r1[34] ;
 wire \rbzero.tex_r1[35] ;
 wire \rbzero.tex_r1[36] ;
 wire \rbzero.tex_r1[37] ;
 wire \rbzero.tex_r1[38] ;
 wire \rbzero.tex_r1[39] ;
 wire \rbzero.tex_r1[3] ;
 wire \rbzero.tex_r1[40] ;
 wire \rbzero.tex_r1[41] ;
 wire \rbzero.tex_r1[42] ;
 wire \rbzero.tex_r1[43] ;
 wire \rbzero.tex_r1[44] ;
 wire \rbzero.tex_r1[45] ;
 wire \rbzero.tex_r1[46] ;
 wire \rbzero.tex_r1[47] ;
 wire \rbzero.tex_r1[48] ;
 wire \rbzero.tex_r1[49] ;
 wire \rbzero.tex_r1[4] ;
 wire \rbzero.tex_r1[50] ;
 wire \rbzero.tex_r1[51] ;
 wire \rbzero.tex_r1[52] ;
 wire \rbzero.tex_r1[53] ;
 wire \rbzero.tex_r1[54] ;
 wire \rbzero.tex_r1[55] ;
 wire \rbzero.tex_r1[56] ;
 wire \rbzero.tex_r1[57] ;
 wire \rbzero.tex_r1[58] ;
 wire \rbzero.tex_r1[59] ;
 wire \rbzero.tex_r1[5] ;
 wire \rbzero.tex_r1[60] ;
 wire \rbzero.tex_r1[61] ;
 wire \rbzero.tex_r1[62] ;
 wire \rbzero.tex_r1[63] ;
 wire \rbzero.tex_r1[6] ;
 wire \rbzero.tex_r1[7] ;
 wire \rbzero.tex_r1[8] ;
 wire \rbzero.tex_r1[9] ;
 wire \rbzero.traced_texVinit[0] ;
 wire \rbzero.traced_texVinit[10] ;
 wire \rbzero.traced_texVinit[11] ;
 wire \rbzero.traced_texVinit[1] ;
 wire \rbzero.traced_texVinit[2] ;
 wire \rbzero.traced_texVinit[3] ;
 wire \rbzero.traced_texVinit[4] ;
 wire \rbzero.traced_texVinit[5] ;
 wire \rbzero.traced_texVinit[6] ;
 wire \rbzero.traced_texVinit[7] ;
 wire \rbzero.traced_texVinit[8] ;
 wire \rbzero.traced_texVinit[9] ;
 wire \rbzero.traced_texa[-10] ;
 wire \rbzero.traced_texa[-11] ;
 wire \rbzero.traced_texa[-12] ;
 wire \rbzero.traced_texa[-1] ;
 wire \rbzero.traced_texa[-2] ;
 wire \rbzero.traced_texa[-3] ;
 wire \rbzero.traced_texa[-4] ;
 wire \rbzero.traced_texa[-5] ;
 wire \rbzero.traced_texa[-6] ;
 wire \rbzero.traced_texa[-7] ;
 wire \rbzero.traced_texa[-8] ;
 wire \rbzero.traced_texa[-9] ;
 wire \rbzero.traced_texa[0] ;
 wire \rbzero.traced_texa[10] ;
 wire \rbzero.traced_texa[11] ;
 wire \rbzero.traced_texa[1] ;
 wire \rbzero.traced_texa[2] ;
 wire \rbzero.traced_texa[3] ;
 wire \rbzero.traced_texa[4] ;
 wire \rbzero.traced_texa[5] ;
 wire \rbzero.traced_texa[6] ;
 wire \rbzero.traced_texa[7] ;
 wire \rbzero.traced_texa[8] ;
 wire \rbzero.traced_texa[9] ;
 wire \rbzero.vga_sync.vsync ;
 wire \rbzero.wall_tracer.rayAddendX[-1] ;
 wire \rbzero.wall_tracer.rayAddendX[-2] ;
 wire \rbzero.wall_tracer.rayAddendX[-3] ;
 wire \rbzero.wall_tracer.rayAddendX[-4] ;
 wire \rbzero.wall_tracer.rayAddendX[-5] ;
 wire \rbzero.wall_tracer.rayAddendX[-6] ;
 wire \rbzero.wall_tracer.rayAddendX[-7] ;
 wire \rbzero.wall_tracer.rayAddendX[-8] ;
 wire \rbzero.wall_tracer.rayAddendX[-9] ;
 wire \rbzero.wall_tracer.rayAddendX[0] ;
 wire \rbzero.wall_tracer.rayAddendX[10] ;
 wire \rbzero.wall_tracer.rayAddendX[11] ;
 wire \rbzero.wall_tracer.rayAddendX[1] ;
 wire \rbzero.wall_tracer.rayAddendX[2] ;
 wire \rbzero.wall_tracer.rayAddendX[3] ;
 wire \rbzero.wall_tracer.rayAddendX[4] ;
 wire \rbzero.wall_tracer.rayAddendX[5] ;
 wire \rbzero.wall_tracer.rayAddendX[6] ;
 wire \rbzero.wall_tracer.rayAddendX[7] ;
 wire \rbzero.wall_tracer.rayAddendX[8] ;
 wire \rbzero.wall_tracer.rayAddendX[9] ;
 wire \rbzero.wall_tracer.rayAddendY[-1] ;
 wire \rbzero.wall_tracer.rayAddendY[-2] ;
 wire \rbzero.wall_tracer.rayAddendY[-3] ;
 wire \rbzero.wall_tracer.rayAddendY[-4] ;
 wire \rbzero.wall_tracer.rayAddendY[-5] ;
 wire \rbzero.wall_tracer.rayAddendY[-6] ;
 wire \rbzero.wall_tracer.rayAddendY[-7] ;
 wire \rbzero.wall_tracer.rayAddendY[-8] ;
 wire \rbzero.wall_tracer.rayAddendY[-9] ;
 wire \rbzero.wall_tracer.rayAddendY[0] ;
 wire \rbzero.wall_tracer.rayAddendY[10] ;
 wire \rbzero.wall_tracer.rayAddendY[11] ;
 wire \rbzero.wall_tracer.rayAddendY[1] ;
 wire \rbzero.wall_tracer.rayAddendY[2] ;
 wire \rbzero.wall_tracer.rayAddendY[3] ;
 wire \rbzero.wall_tracer.rayAddendY[4] ;
 wire \rbzero.wall_tracer.rayAddendY[5] ;
 wire \rbzero.wall_tracer.rayAddendY[6] ;
 wire \rbzero.wall_tracer.rayAddendY[7] ;
 wire \rbzero.wall_tracer.rayAddendY[8] ;
 wire \rbzero.wall_tracer.rayAddendY[9] ;
 wire \rbzero.wall_tracer.rcp_sel[0] ;
 wire \rbzero.wall_tracer.rcp_sel[2] ;
 wire \rbzero.wall_tracer.side ;
 wire \rbzero.wall_tracer.state[0] ;
 wire \rbzero.wall_tracer.state[10] ;
 wire \rbzero.wall_tracer.state[11] ;
 wire \rbzero.wall_tracer.state[12] ;
 wire \rbzero.wall_tracer.state[13] ;
 wire \rbzero.wall_tracer.state[14] ;
 wire \rbzero.wall_tracer.state[1] ;
 wire \rbzero.wall_tracer.state[2] ;
 wire \rbzero.wall_tracer.state[3] ;
 wire \rbzero.wall_tracer.state[4] ;
 wire \rbzero.wall_tracer.state[5] ;
 wire \rbzero.wall_tracer.state[6] ;
 wire \rbzero.wall_tracer.state[7] ;
 wire \rbzero.wall_tracer.state[8] ;
 wire \rbzero.wall_tracer.state[9] ;
 wire \rbzero.wall_tracer.stepDistX[-10] ;
 wire \rbzero.wall_tracer.stepDistX[-11] ;
 wire \rbzero.wall_tracer.stepDistX[-12] ;
 wire \rbzero.wall_tracer.stepDistX[-1] ;
 wire \rbzero.wall_tracer.stepDistX[-2] ;
 wire \rbzero.wall_tracer.stepDistX[-3] ;
 wire \rbzero.wall_tracer.stepDistX[-4] ;
 wire \rbzero.wall_tracer.stepDistX[-5] ;
 wire \rbzero.wall_tracer.stepDistX[-6] ;
 wire \rbzero.wall_tracer.stepDistX[-7] ;
 wire \rbzero.wall_tracer.stepDistX[-8] ;
 wire \rbzero.wall_tracer.stepDistX[-9] ;
 wire \rbzero.wall_tracer.stepDistX[0] ;
 wire \rbzero.wall_tracer.stepDistX[10] ;
 wire \rbzero.wall_tracer.stepDistX[11] ;
 wire \rbzero.wall_tracer.stepDistX[1] ;
 wire \rbzero.wall_tracer.stepDistX[2] ;
 wire \rbzero.wall_tracer.stepDistX[3] ;
 wire \rbzero.wall_tracer.stepDistX[4] ;
 wire \rbzero.wall_tracer.stepDistX[5] ;
 wire \rbzero.wall_tracer.stepDistX[6] ;
 wire \rbzero.wall_tracer.stepDistX[7] ;
 wire \rbzero.wall_tracer.stepDistX[8] ;
 wire \rbzero.wall_tracer.stepDistX[9] ;
 wire \rbzero.wall_tracer.stepDistY[-10] ;
 wire \rbzero.wall_tracer.stepDistY[-11] ;
 wire \rbzero.wall_tracer.stepDistY[-12] ;
 wire \rbzero.wall_tracer.stepDistY[-1] ;
 wire \rbzero.wall_tracer.stepDistY[-2] ;
 wire \rbzero.wall_tracer.stepDistY[-3] ;
 wire \rbzero.wall_tracer.stepDistY[-4] ;
 wire \rbzero.wall_tracer.stepDistY[-5] ;
 wire \rbzero.wall_tracer.stepDistY[-6] ;
 wire \rbzero.wall_tracer.stepDistY[-7] ;
 wire \rbzero.wall_tracer.stepDistY[-8] ;
 wire \rbzero.wall_tracer.stepDistY[-9] ;
 wire \rbzero.wall_tracer.stepDistY[0] ;
 wire \rbzero.wall_tracer.stepDistY[10] ;
 wire \rbzero.wall_tracer.stepDistY[11] ;
 wire \rbzero.wall_tracer.stepDistY[1] ;
 wire \rbzero.wall_tracer.stepDistY[2] ;
 wire \rbzero.wall_tracer.stepDistY[3] ;
 wire \rbzero.wall_tracer.stepDistY[4] ;
 wire \rbzero.wall_tracer.stepDistY[5] ;
 wire \rbzero.wall_tracer.stepDistY[6] ;
 wire \rbzero.wall_tracer.stepDistY[7] ;
 wire \rbzero.wall_tracer.stepDistY[8] ;
 wire \rbzero.wall_tracer.stepDistY[9] ;
 wire \rbzero.wall_tracer.texu[0] ;
 wire \rbzero.wall_tracer.texu[1] ;
 wire \rbzero.wall_tracer.texu[2] ;
 wire \rbzero.wall_tracer.texu[3] ;
 wire \rbzero.wall_tracer.texu[4] ;
 wire \rbzero.wall_tracer.texu[5] ;
 wire \rbzero.wall_tracer.trackDistX[-10] ;
 wire \rbzero.wall_tracer.trackDistX[-11] ;
 wire \rbzero.wall_tracer.trackDistX[-12] ;
 wire \rbzero.wall_tracer.trackDistX[-1] ;
 wire \rbzero.wall_tracer.trackDistX[-2] ;
 wire \rbzero.wall_tracer.trackDistX[-3] ;
 wire \rbzero.wall_tracer.trackDistX[-4] ;
 wire \rbzero.wall_tracer.trackDistX[-5] ;
 wire \rbzero.wall_tracer.trackDistX[-6] ;
 wire \rbzero.wall_tracer.trackDistX[-7] ;
 wire \rbzero.wall_tracer.trackDistX[-8] ;
 wire \rbzero.wall_tracer.trackDistX[-9] ;
 wire \rbzero.wall_tracer.trackDistX[0] ;
 wire \rbzero.wall_tracer.trackDistX[10] ;
 wire \rbzero.wall_tracer.trackDistX[11] ;
 wire \rbzero.wall_tracer.trackDistX[1] ;
 wire \rbzero.wall_tracer.trackDistX[2] ;
 wire \rbzero.wall_tracer.trackDistX[3] ;
 wire \rbzero.wall_tracer.trackDistX[4] ;
 wire \rbzero.wall_tracer.trackDistX[5] ;
 wire \rbzero.wall_tracer.trackDistX[6] ;
 wire \rbzero.wall_tracer.trackDistX[7] ;
 wire \rbzero.wall_tracer.trackDistX[8] ;
 wire \rbzero.wall_tracer.trackDistX[9] ;
 wire \rbzero.wall_tracer.trackDistY[-10] ;
 wire \rbzero.wall_tracer.trackDistY[-11] ;
 wire \rbzero.wall_tracer.trackDistY[-12] ;
 wire \rbzero.wall_tracer.trackDistY[-1] ;
 wire \rbzero.wall_tracer.trackDistY[-2] ;
 wire \rbzero.wall_tracer.trackDistY[-3] ;
 wire \rbzero.wall_tracer.trackDistY[-4] ;
 wire \rbzero.wall_tracer.trackDistY[-5] ;
 wire \rbzero.wall_tracer.trackDistY[-6] ;
 wire \rbzero.wall_tracer.trackDistY[-7] ;
 wire \rbzero.wall_tracer.trackDistY[-8] ;
 wire \rbzero.wall_tracer.trackDistY[-9] ;
 wire \rbzero.wall_tracer.trackDistY[0] ;
 wire \rbzero.wall_tracer.trackDistY[10] ;
 wire \rbzero.wall_tracer.trackDistY[11] ;
 wire \rbzero.wall_tracer.trackDistY[1] ;
 wire \rbzero.wall_tracer.trackDistY[2] ;
 wire \rbzero.wall_tracer.trackDistY[3] ;
 wire \rbzero.wall_tracer.trackDistY[4] ;
 wire \rbzero.wall_tracer.trackDistY[5] ;
 wire \rbzero.wall_tracer.trackDistY[6] ;
 wire \rbzero.wall_tracer.trackDistY[7] ;
 wire \rbzero.wall_tracer.trackDistY[8] ;
 wire \rbzero.wall_tracer.trackDistY[9] ;
 wire \rbzero.wall_tracer.visualWallDist[-10] ;
 wire \rbzero.wall_tracer.visualWallDist[-11] ;
 wire \rbzero.wall_tracer.visualWallDist[-12] ;
 wire \rbzero.wall_tracer.visualWallDist[-1] ;
 wire \rbzero.wall_tracer.visualWallDist[-2] ;
 wire \rbzero.wall_tracer.visualWallDist[-3] ;
 wire \rbzero.wall_tracer.visualWallDist[-4] ;
 wire \rbzero.wall_tracer.visualWallDist[-5] ;
 wire \rbzero.wall_tracer.visualWallDist[-6] ;
 wire \rbzero.wall_tracer.visualWallDist[-7] ;
 wire \rbzero.wall_tracer.visualWallDist[-8] ;
 wire \rbzero.wall_tracer.visualWallDist[-9] ;
 wire \rbzero.wall_tracer.visualWallDist[0] ;
 wire \rbzero.wall_tracer.visualWallDist[10] ;
 wire \rbzero.wall_tracer.visualWallDist[11] ;
 wire \rbzero.wall_tracer.visualWallDist[1] ;
 wire \rbzero.wall_tracer.visualWallDist[2] ;
 wire \rbzero.wall_tracer.visualWallDist[3] ;
 wire \rbzero.wall_tracer.visualWallDist[4] ;
 wire \rbzero.wall_tracer.visualWallDist[5] ;
 wire \rbzero.wall_tracer.visualWallDist[6] ;
 wire \rbzero.wall_tracer.visualWallDist[7] ;
 wire \rbzero.wall_tracer.visualWallDist[8] ;
 wire \rbzero.wall_tracer.visualWallDist[9] ;
 wire \rbzero.wall_tracer.wall[0] ;
 wire \rbzero.wall_tracer.wall[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;

 sky130_fd_sc_hd__clkbuf_4 _10175_ (.A(\gpout0.hpos[0] ),
    .X(_03288_));
 sky130_fd_sc_hd__clkbuf_2 _10176_ (.A(_03288_),
    .X(_03289_));
 sky130_fd_sc_hd__clkbuf_4 _10177_ (.A(\gpout0.hpos[7] ),
    .X(_03290_));
 sky130_fd_sc_hd__clkbuf_4 _10178_ (.A(_03290_),
    .X(_03291_));
 sky130_fd_sc_hd__xor2_4 _10179_ (.A(net46),
    .B(net45),
    .X(_03292_));
 sky130_fd_sc_hd__clkbuf_4 _10180_ (.A(\gpout0.hpos[8] ),
    .X(_03293_));
 sky130_fd_sc_hd__buf_2 _10181_ (.A(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__buf_2 _10182_ (.A(\gpout0.hpos[9] ),
    .X(_03295_));
 sky130_fd_sc_hd__inv_2 _10183_ (.A(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hd__nor2_1 _10184_ (.A(_03294_),
    .B(_03296_),
    .Y(_03297_));
 sky130_fd_sc_hd__and4_2 _10185_ (.A(_03289_),
    .B(_03291_),
    .C(_03292_),
    .D(_03297_),
    .X(_03298_));
 sky130_fd_sc_hd__clkbuf_4 _10186_ (.A(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__clkbuf_4 _10187_ (.A(_03299_),
    .X(_03300_));
 sky130_fd_sc_hd__mux2_1 _10188_ (.A0(\rbzero.tex_b1[63] ),
    .A1(net50),
    .S(_03300_),
    .X(_03301_));
 sky130_fd_sc_hd__clkbuf_1 _10189_ (.A(_03301_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _10190_ (.A0(\rbzero.tex_b1[62] ),
    .A1(\rbzero.tex_b1[63] ),
    .S(_03300_),
    .X(_03302_));
 sky130_fd_sc_hd__clkbuf_1 _10191_ (.A(_03302_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _10192_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[62] ),
    .S(_03300_),
    .X(_03303_));
 sky130_fd_sc_hd__clkbuf_1 _10193_ (.A(_03303_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _10194_ (.A0(\rbzero.tex_b1[60] ),
    .A1(\rbzero.tex_b1[61] ),
    .S(_03300_),
    .X(_03304_));
 sky130_fd_sc_hd__clkbuf_1 _10195_ (.A(_03304_),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _10196_ (.A0(\rbzero.tex_b1[59] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_03300_),
    .X(_03305_));
 sky130_fd_sc_hd__clkbuf_1 _10197_ (.A(_03305_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _10198_ (.A0(\rbzero.tex_b1[58] ),
    .A1(\rbzero.tex_b1[59] ),
    .S(_03300_),
    .X(_03306_));
 sky130_fd_sc_hd__clkbuf_1 _10199_ (.A(_03306_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _10200_ (.A0(\rbzero.tex_b1[57] ),
    .A1(\rbzero.tex_b1[58] ),
    .S(_03300_),
    .X(_03307_));
 sky130_fd_sc_hd__clkbuf_1 _10201_ (.A(_03307_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _10202_ (.A0(\rbzero.tex_b1[56] ),
    .A1(\rbzero.tex_b1[57] ),
    .S(_03300_),
    .X(_03308_));
 sky130_fd_sc_hd__clkbuf_1 _10203_ (.A(_03308_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _10204_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[56] ),
    .S(_03300_),
    .X(_03309_));
 sky130_fd_sc_hd__clkbuf_1 _10205_ (.A(_03309_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _10206_ (.A0(\rbzero.tex_b1[54] ),
    .A1(\rbzero.tex_b1[55] ),
    .S(_03300_),
    .X(_03310_));
 sky130_fd_sc_hd__clkbuf_1 _10207_ (.A(_03310_),
    .X(_01384_));
 sky130_fd_sc_hd__clkbuf_4 _10208_ (.A(_03299_),
    .X(_03311_));
 sky130_fd_sc_hd__mux2_1 _10209_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(_03311_),
    .X(_03312_));
 sky130_fd_sc_hd__clkbuf_1 _10210_ (.A(_03312_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _10211_ (.A0(\rbzero.tex_b1[52] ),
    .A1(\rbzero.tex_b1[53] ),
    .S(_03311_),
    .X(_03313_));
 sky130_fd_sc_hd__clkbuf_1 _10212_ (.A(_03313_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _10213_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(_03311_),
    .X(_03314_));
 sky130_fd_sc_hd__clkbuf_1 _10214_ (.A(_03314_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _10215_ (.A0(\rbzero.tex_b1[50] ),
    .A1(\rbzero.tex_b1[51] ),
    .S(_03311_),
    .X(_03315_));
 sky130_fd_sc_hd__clkbuf_1 _10216_ (.A(_03315_),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _10217_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_03311_),
    .X(_03316_));
 sky130_fd_sc_hd__clkbuf_1 _10218_ (.A(_03316_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _10219_ (.A0(\rbzero.tex_b1[48] ),
    .A1(\rbzero.tex_b1[49] ),
    .S(_03311_),
    .X(_03317_));
 sky130_fd_sc_hd__clkbuf_1 _10220_ (.A(_03317_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _10221_ (.A0(\rbzero.tex_b1[47] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(_03311_),
    .X(_03318_));
 sky130_fd_sc_hd__clkbuf_1 _10222_ (.A(_03318_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _10223_ (.A0(\rbzero.tex_b1[46] ),
    .A1(\rbzero.tex_b1[47] ),
    .S(_03311_),
    .X(_03319_));
 sky130_fd_sc_hd__clkbuf_1 _10224_ (.A(_03319_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _10225_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[46] ),
    .S(_03311_),
    .X(_03320_));
 sky130_fd_sc_hd__clkbuf_1 _10226_ (.A(_03320_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _10227_ (.A0(\rbzero.tex_b1[44] ),
    .A1(\rbzero.tex_b1[45] ),
    .S(_03311_),
    .X(_03321_));
 sky130_fd_sc_hd__clkbuf_1 _10228_ (.A(_03321_),
    .X(_01374_));
 sky130_fd_sc_hd__clkbuf_4 _10229_ (.A(_03299_),
    .X(_03322_));
 sky130_fd_sc_hd__mux2_1 _10230_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__clkbuf_1 _10231_ (.A(_03323_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _10232_ (.A0(\rbzero.tex_b1[42] ),
    .A1(\rbzero.tex_b1[43] ),
    .S(_03322_),
    .X(_03324_));
 sky130_fd_sc_hd__clkbuf_1 _10233_ (.A(_03324_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _10234_ (.A0(\rbzero.tex_b1[41] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(_03322_),
    .X(_03325_));
 sky130_fd_sc_hd__clkbuf_1 _10235_ (.A(_03325_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _10236_ (.A0(\rbzero.tex_b1[40] ),
    .A1(\rbzero.tex_b1[41] ),
    .S(_03322_),
    .X(_03326_));
 sky130_fd_sc_hd__clkbuf_1 _10237_ (.A(_03326_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _10238_ (.A0(\rbzero.tex_b1[39] ),
    .A1(\rbzero.tex_b1[40] ),
    .S(_03322_),
    .X(_03327_));
 sky130_fd_sc_hd__clkbuf_1 _10239_ (.A(_03327_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _10240_ (.A0(\rbzero.tex_b1[38] ),
    .A1(\rbzero.tex_b1[39] ),
    .S(_03322_),
    .X(_03328_));
 sky130_fd_sc_hd__clkbuf_1 _10241_ (.A(_03328_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _10242_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[38] ),
    .S(_03322_),
    .X(_03329_));
 sky130_fd_sc_hd__clkbuf_1 _10243_ (.A(_03329_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _10244_ (.A0(\rbzero.tex_b1[36] ),
    .A1(\rbzero.tex_b1[37] ),
    .S(_03322_),
    .X(_03330_));
 sky130_fd_sc_hd__clkbuf_1 _10245_ (.A(_03330_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _10246_ (.A0(\rbzero.tex_b1[35] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(_03322_),
    .X(_03331_));
 sky130_fd_sc_hd__clkbuf_1 _10247_ (.A(_03331_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _10248_ (.A0(\rbzero.tex_b1[34] ),
    .A1(\rbzero.tex_b1[35] ),
    .S(_03322_),
    .X(_03332_));
 sky130_fd_sc_hd__clkbuf_1 _10249_ (.A(_03332_),
    .X(_01364_));
 sky130_fd_sc_hd__clkbuf_4 _10250_ (.A(_03299_),
    .X(_03333_));
 sky130_fd_sc_hd__mux2_1 _10251_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[34] ),
    .S(_03333_),
    .X(_03334_));
 sky130_fd_sc_hd__clkbuf_1 _10252_ (.A(_03334_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _10253_ (.A0(\rbzero.tex_b1[32] ),
    .A1(\rbzero.tex_b1[33] ),
    .S(_03333_),
    .X(_03335_));
 sky130_fd_sc_hd__clkbuf_1 _10254_ (.A(_03335_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _10255_ (.A0(\rbzero.tex_b1[31] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(_03333_),
    .X(_03336_));
 sky130_fd_sc_hd__clkbuf_1 _10256_ (.A(_03336_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _10257_ (.A0(\rbzero.tex_b1[30] ),
    .A1(\rbzero.tex_b1[31] ),
    .S(_03333_),
    .X(_03337_));
 sky130_fd_sc_hd__clkbuf_1 _10258_ (.A(_03337_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _10259_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[30] ),
    .S(_03333_),
    .X(_03338_));
 sky130_fd_sc_hd__clkbuf_1 _10260_ (.A(_03338_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _10261_ (.A0(\rbzero.tex_b1[28] ),
    .A1(\rbzero.tex_b1[29] ),
    .S(_03333_),
    .X(_03339_));
 sky130_fd_sc_hd__clkbuf_1 _10262_ (.A(_03339_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _10263_ (.A0(\rbzero.tex_b1[27] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(_03333_),
    .X(_03340_));
 sky130_fd_sc_hd__clkbuf_1 _10264_ (.A(_03340_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _10265_ (.A0(\rbzero.tex_b1[26] ),
    .A1(\rbzero.tex_b1[27] ),
    .S(_03333_),
    .X(_03341_));
 sky130_fd_sc_hd__clkbuf_1 _10266_ (.A(_03341_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _10267_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[26] ),
    .S(_03333_),
    .X(_03342_));
 sky130_fd_sc_hd__clkbuf_1 _10268_ (.A(_03342_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _10269_ (.A0(\rbzero.tex_b1[24] ),
    .A1(\rbzero.tex_b1[25] ),
    .S(_03333_),
    .X(_03343_));
 sky130_fd_sc_hd__clkbuf_1 _10270_ (.A(_03343_),
    .X(_01354_));
 sky130_fd_sc_hd__clkbuf_4 _10271_ (.A(_03299_),
    .X(_03344_));
 sky130_fd_sc_hd__mux2_1 _10272_ (.A0(\rbzero.tex_b1[23] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(_03344_),
    .X(_03345_));
 sky130_fd_sc_hd__clkbuf_1 _10273_ (.A(_03345_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _10274_ (.A0(\rbzero.tex_b1[22] ),
    .A1(\rbzero.tex_b1[23] ),
    .S(_03344_),
    .X(_03346_));
 sky130_fd_sc_hd__clkbuf_1 _10275_ (.A(_03346_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _10276_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[22] ),
    .S(_03344_),
    .X(_03347_));
 sky130_fd_sc_hd__clkbuf_1 _10277_ (.A(_03347_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _10278_ (.A0(\rbzero.tex_b1[20] ),
    .A1(\rbzero.tex_b1[21] ),
    .S(_03344_),
    .X(_03348_));
 sky130_fd_sc_hd__clkbuf_1 _10279_ (.A(_03348_),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _10280_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(_03344_),
    .X(_03349_));
 sky130_fd_sc_hd__clkbuf_1 _10281_ (.A(_03349_),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _10282_ (.A0(\rbzero.tex_b1[18] ),
    .A1(\rbzero.tex_b1[19] ),
    .S(_03344_),
    .X(_03350_));
 sky130_fd_sc_hd__clkbuf_1 _10283_ (.A(_03350_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _10284_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(_03344_),
    .X(_03351_));
 sky130_fd_sc_hd__clkbuf_1 _10285_ (.A(_03351_),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _10286_ (.A0(\rbzero.tex_b1[16] ),
    .A1(\rbzero.tex_b1[17] ),
    .S(_03344_),
    .X(_03352_));
 sky130_fd_sc_hd__clkbuf_1 _10287_ (.A(_03352_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _10288_ (.A0(\rbzero.tex_b1[15] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(_03344_),
    .X(_03353_));
 sky130_fd_sc_hd__clkbuf_1 _10289_ (.A(_03353_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _10290_ (.A0(\rbzero.tex_b1[14] ),
    .A1(\rbzero.tex_b1[15] ),
    .S(_03344_),
    .X(_03354_));
 sky130_fd_sc_hd__clkbuf_1 _10291_ (.A(_03354_),
    .X(_01344_));
 sky130_fd_sc_hd__clkbuf_4 _10292_ (.A(_03299_),
    .X(_03355_));
 sky130_fd_sc_hd__mux2_1 _10293_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[14] ),
    .S(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__clkbuf_1 _10294_ (.A(_03356_),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _10295_ (.A0(\rbzero.tex_b1[12] ),
    .A1(\rbzero.tex_b1[13] ),
    .S(_03355_),
    .X(_03357_));
 sky130_fd_sc_hd__clkbuf_1 _10296_ (.A(_03357_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _10297_ (.A0(\rbzero.tex_b1[11] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_03355_),
    .X(_03358_));
 sky130_fd_sc_hd__clkbuf_1 _10298_ (.A(_03358_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _10299_ (.A0(\rbzero.tex_b1[10] ),
    .A1(\rbzero.tex_b1[11] ),
    .S(_03355_),
    .X(_03359_));
 sky130_fd_sc_hd__clkbuf_1 _10300_ (.A(_03359_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _10301_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[10] ),
    .S(_03355_),
    .X(_03360_));
 sky130_fd_sc_hd__clkbuf_1 _10302_ (.A(_03360_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _10303_ (.A0(\rbzero.tex_b1[8] ),
    .A1(\rbzero.tex_b1[9] ),
    .S(_03355_),
    .X(_03361_));
 sky130_fd_sc_hd__clkbuf_1 _10304_ (.A(_03361_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _10305_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_03355_),
    .X(_03362_));
 sky130_fd_sc_hd__clkbuf_1 _10306_ (.A(_03362_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _10307_ (.A0(\rbzero.tex_b1[6] ),
    .A1(\rbzero.tex_b1[7] ),
    .S(_03355_),
    .X(_03363_));
 sky130_fd_sc_hd__clkbuf_1 _10308_ (.A(_03363_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _10309_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(_03355_),
    .X(_03364_));
 sky130_fd_sc_hd__clkbuf_1 _10310_ (.A(_03364_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _10311_ (.A0(\rbzero.tex_b1[4] ),
    .A1(\rbzero.tex_b1[5] ),
    .S(_03355_),
    .X(_03365_));
 sky130_fd_sc_hd__clkbuf_1 _10312_ (.A(_03365_),
    .X(_01334_));
 sky130_fd_sc_hd__clkbuf_4 _10313_ (.A(_03299_),
    .X(_03366_));
 sky130_fd_sc_hd__mux2_1 _10314_ (.A0(\rbzero.tex_b1[3] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_03366_),
    .X(_03367_));
 sky130_fd_sc_hd__clkbuf_1 _10315_ (.A(_03367_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _10316_ (.A0(\rbzero.tex_b1[2] ),
    .A1(\rbzero.tex_b1[3] ),
    .S(_03366_),
    .X(_03368_));
 sky130_fd_sc_hd__clkbuf_1 _10317_ (.A(_03368_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _10318_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[2] ),
    .S(_03366_),
    .X(_03369_));
 sky130_fd_sc_hd__clkbuf_1 _10319_ (.A(_03369_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _10320_ (.A0(\rbzero.tex_b1[0] ),
    .A1(\rbzero.tex_b1[1] ),
    .S(_03366_),
    .X(_03370_));
 sky130_fd_sc_hd__clkbuf_1 _10321_ (.A(_03370_),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _10322_ (.A0(\rbzero.tex_r1[63] ),
    .A1(net48),
    .S(_03366_),
    .X(_03371_));
 sky130_fd_sc_hd__clkbuf_1 _10323_ (.A(_03371_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _10324_ (.A0(\rbzero.tex_r1[62] ),
    .A1(\rbzero.tex_r1[63] ),
    .S(_03366_),
    .X(_03372_));
 sky130_fd_sc_hd__clkbuf_1 _10325_ (.A(_03372_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _10326_ (.A0(\rbzero.tex_r1[61] ),
    .A1(\rbzero.tex_r1[62] ),
    .S(_03366_),
    .X(_03373_));
 sky130_fd_sc_hd__clkbuf_1 _10327_ (.A(_03373_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _10328_ (.A0(\rbzero.tex_r1[60] ),
    .A1(\rbzero.tex_r1[61] ),
    .S(_03366_),
    .X(_03374_));
 sky130_fd_sc_hd__clkbuf_1 _10329_ (.A(_03374_),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _10330_ (.A0(\rbzero.tex_r1[59] ),
    .A1(\rbzero.tex_r1[60] ),
    .S(_03366_),
    .X(_03375_));
 sky130_fd_sc_hd__clkbuf_1 _10331_ (.A(_03375_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _10332_ (.A0(\rbzero.tex_r1[58] ),
    .A1(\rbzero.tex_r1[59] ),
    .S(_03366_),
    .X(_03376_));
 sky130_fd_sc_hd__clkbuf_1 _10333_ (.A(_03376_),
    .X(_01298_));
 sky130_fd_sc_hd__clkbuf_4 _10334_ (.A(_03299_),
    .X(_03377_));
 sky130_fd_sc_hd__mux2_1 _10335_ (.A0(\rbzero.tex_r1[57] ),
    .A1(\rbzero.tex_r1[58] ),
    .S(_03377_),
    .X(_03378_));
 sky130_fd_sc_hd__clkbuf_1 _10336_ (.A(_03378_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _10337_ (.A0(\rbzero.tex_r1[56] ),
    .A1(\rbzero.tex_r1[57] ),
    .S(_03377_),
    .X(_03379_));
 sky130_fd_sc_hd__clkbuf_1 _10338_ (.A(_03379_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _10339_ (.A0(\rbzero.tex_r1[55] ),
    .A1(\rbzero.tex_r1[56] ),
    .S(_03377_),
    .X(_03380_));
 sky130_fd_sc_hd__clkbuf_1 _10340_ (.A(_03380_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _10341_ (.A0(\rbzero.tex_r1[54] ),
    .A1(\rbzero.tex_r1[55] ),
    .S(_03377_),
    .X(_03381_));
 sky130_fd_sc_hd__clkbuf_1 _10342_ (.A(_03381_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _10343_ (.A0(\rbzero.tex_r1[53] ),
    .A1(\rbzero.tex_r1[54] ),
    .S(_03377_),
    .X(_03382_));
 sky130_fd_sc_hd__clkbuf_1 _10344_ (.A(_03382_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _10345_ (.A0(\rbzero.tex_r1[52] ),
    .A1(\rbzero.tex_r1[53] ),
    .S(_03377_),
    .X(_03383_));
 sky130_fd_sc_hd__clkbuf_1 _10346_ (.A(_03383_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _10347_ (.A0(\rbzero.tex_r1[51] ),
    .A1(\rbzero.tex_r1[52] ),
    .S(_03377_),
    .X(_03384_));
 sky130_fd_sc_hd__clkbuf_1 _10348_ (.A(_03384_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _10349_ (.A0(\rbzero.tex_r1[50] ),
    .A1(\rbzero.tex_r1[51] ),
    .S(_03377_),
    .X(_03385_));
 sky130_fd_sc_hd__clkbuf_1 _10350_ (.A(_03385_),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _10351_ (.A0(\rbzero.tex_r1[49] ),
    .A1(\rbzero.tex_r1[50] ),
    .S(_03377_),
    .X(_03386_));
 sky130_fd_sc_hd__clkbuf_1 _10352_ (.A(_03386_),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _10353_ (.A0(\rbzero.tex_r1[48] ),
    .A1(\rbzero.tex_r1[49] ),
    .S(_03377_),
    .X(_03387_));
 sky130_fd_sc_hd__clkbuf_1 _10354_ (.A(_03387_),
    .X(_01288_));
 sky130_fd_sc_hd__clkbuf_4 _10355_ (.A(_03298_),
    .X(_03388_));
 sky130_fd_sc_hd__clkbuf_4 _10356_ (.A(_03388_),
    .X(_03389_));
 sky130_fd_sc_hd__mux2_1 _10357_ (.A0(\rbzero.tex_r1[47] ),
    .A1(\rbzero.tex_r1[48] ),
    .S(_03389_),
    .X(_03390_));
 sky130_fd_sc_hd__clkbuf_1 _10358_ (.A(_03390_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _10359_ (.A0(\rbzero.tex_r1[46] ),
    .A1(\rbzero.tex_r1[47] ),
    .S(_03389_),
    .X(_03391_));
 sky130_fd_sc_hd__clkbuf_1 _10360_ (.A(_03391_),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _10361_ (.A0(\rbzero.tex_r1[45] ),
    .A1(\rbzero.tex_r1[46] ),
    .S(_03389_),
    .X(_03392_));
 sky130_fd_sc_hd__clkbuf_1 _10362_ (.A(_03392_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _10363_ (.A0(\rbzero.tex_r1[44] ),
    .A1(\rbzero.tex_r1[45] ),
    .S(_03389_),
    .X(_03393_));
 sky130_fd_sc_hd__clkbuf_1 _10364_ (.A(_03393_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _10365_ (.A0(\rbzero.tex_r1[43] ),
    .A1(\rbzero.tex_r1[44] ),
    .S(_03389_),
    .X(_03394_));
 sky130_fd_sc_hd__clkbuf_1 _10366_ (.A(_03394_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _10367_ (.A0(\rbzero.tex_r1[42] ),
    .A1(\rbzero.tex_r1[43] ),
    .S(_03389_),
    .X(_03395_));
 sky130_fd_sc_hd__clkbuf_1 _10368_ (.A(_03395_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _10369_ (.A0(\rbzero.tex_r1[41] ),
    .A1(\rbzero.tex_r1[42] ),
    .S(_03389_),
    .X(_03396_));
 sky130_fd_sc_hd__clkbuf_1 _10370_ (.A(_03396_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _10371_ (.A0(\rbzero.tex_r1[40] ),
    .A1(\rbzero.tex_r1[41] ),
    .S(_03389_),
    .X(_03397_));
 sky130_fd_sc_hd__clkbuf_1 _10372_ (.A(_03397_),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _10373_ (.A0(\rbzero.tex_r1[39] ),
    .A1(\rbzero.tex_r1[40] ),
    .S(_03389_),
    .X(_03398_));
 sky130_fd_sc_hd__clkbuf_1 _10374_ (.A(_03398_),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _10375_ (.A0(\rbzero.tex_r1[38] ),
    .A1(\rbzero.tex_r1[39] ),
    .S(_03389_),
    .X(_03399_));
 sky130_fd_sc_hd__clkbuf_1 _10376_ (.A(_03399_),
    .X(_01278_));
 sky130_fd_sc_hd__clkbuf_4 _10377_ (.A(_03388_),
    .X(_03400_));
 sky130_fd_sc_hd__mux2_1 _10378_ (.A0(\rbzero.tex_r1[37] ),
    .A1(\rbzero.tex_r1[38] ),
    .S(_03400_),
    .X(_03401_));
 sky130_fd_sc_hd__clkbuf_1 _10379_ (.A(_03401_),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _10380_ (.A0(\rbzero.tex_r1[36] ),
    .A1(\rbzero.tex_r1[37] ),
    .S(_03400_),
    .X(_03402_));
 sky130_fd_sc_hd__clkbuf_1 _10381_ (.A(_03402_),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _10382_ (.A0(\rbzero.tex_r1[35] ),
    .A1(\rbzero.tex_r1[36] ),
    .S(_03400_),
    .X(_03403_));
 sky130_fd_sc_hd__clkbuf_1 _10383_ (.A(_03403_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _10384_ (.A0(\rbzero.tex_r1[34] ),
    .A1(\rbzero.tex_r1[35] ),
    .S(_03400_),
    .X(_03404_));
 sky130_fd_sc_hd__clkbuf_1 _10385_ (.A(_03404_),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _10386_ (.A0(\rbzero.tex_r1[33] ),
    .A1(\rbzero.tex_r1[34] ),
    .S(_03400_),
    .X(_03405_));
 sky130_fd_sc_hd__clkbuf_1 _10387_ (.A(_03405_),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _10388_ (.A0(\rbzero.tex_r1[32] ),
    .A1(\rbzero.tex_r1[33] ),
    .S(_03400_),
    .X(_03406_));
 sky130_fd_sc_hd__clkbuf_1 _10389_ (.A(_03406_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _10390_ (.A0(\rbzero.tex_r1[31] ),
    .A1(\rbzero.tex_r1[32] ),
    .S(_03400_),
    .X(_03407_));
 sky130_fd_sc_hd__clkbuf_1 _10391_ (.A(_03407_),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _10392_ (.A0(\rbzero.tex_r1[30] ),
    .A1(\rbzero.tex_r1[31] ),
    .S(_03400_),
    .X(_03408_));
 sky130_fd_sc_hd__clkbuf_1 _10393_ (.A(_03408_),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _10394_ (.A0(\rbzero.tex_r1[29] ),
    .A1(\rbzero.tex_r1[30] ),
    .S(_03400_),
    .X(_03409_));
 sky130_fd_sc_hd__clkbuf_1 _10395_ (.A(_03409_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _10396_ (.A0(\rbzero.tex_r1[28] ),
    .A1(\rbzero.tex_r1[29] ),
    .S(_03400_),
    .X(_03410_));
 sky130_fd_sc_hd__clkbuf_1 _10397_ (.A(_03410_),
    .X(_01268_));
 sky130_fd_sc_hd__clkbuf_4 _10398_ (.A(_03388_),
    .X(_03411_));
 sky130_fd_sc_hd__mux2_1 _10399_ (.A0(\rbzero.tex_r1[27] ),
    .A1(\rbzero.tex_r1[28] ),
    .S(_03411_),
    .X(_03412_));
 sky130_fd_sc_hd__clkbuf_1 _10400_ (.A(_03412_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _10401_ (.A0(\rbzero.tex_r1[26] ),
    .A1(\rbzero.tex_r1[27] ),
    .S(_03411_),
    .X(_03413_));
 sky130_fd_sc_hd__clkbuf_1 _10402_ (.A(_03413_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _10403_ (.A0(\rbzero.tex_r1[25] ),
    .A1(\rbzero.tex_r1[26] ),
    .S(_03411_),
    .X(_03414_));
 sky130_fd_sc_hd__clkbuf_1 _10404_ (.A(_03414_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _10405_ (.A0(\rbzero.tex_r1[24] ),
    .A1(\rbzero.tex_r1[25] ),
    .S(_03411_),
    .X(_03415_));
 sky130_fd_sc_hd__clkbuf_1 _10406_ (.A(_03415_),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _10407_ (.A0(\rbzero.tex_r1[23] ),
    .A1(\rbzero.tex_r1[24] ),
    .S(_03411_),
    .X(_03416_));
 sky130_fd_sc_hd__clkbuf_1 _10408_ (.A(_03416_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _10409_ (.A0(\rbzero.tex_r1[22] ),
    .A1(\rbzero.tex_r1[23] ),
    .S(_03411_),
    .X(_03417_));
 sky130_fd_sc_hd__clkbuf_1 _10410_ (.A(_03417_),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_1 _10411_ (.A0(\rbzero.tex_r1[21] ),
    .A1(\rbzero.tex_r1[22] ),
    .S(_03411_),
    .X(_03418_));
 sky130_fd_sc_hd__clkbuf_1 _10412_ (.A(_03418_),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _10413_ (.A0(\rbzero.tex_r1[20] ),
    .A1(\rbzero.tex_r1[21] ),
    .S(_03411_),
    .X(_03419_));
 sky130_fd_sc_hd__clkbuf_1 _10414_ (.A(_03419_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _10415_ (.A0(\rbzero.tex_r1[19] ),
    .A1(\rbzero.tex_r1[20] ),
    .S(_03411_),
    .X(_03420_));
 sky130_fd_sc_hd__clkbuf_1 _10416_ (.A(_03420_),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _10417_ (.A0(\rbzero.tex_r1[18] ),
    .A1(\rbzero.tex_r1[19] ),
    .S(_03411_),
    .X(_03421_));
 sky130_fd_sc_hd__clkbuf_1 _10418_ (.A(_03421_),
    .X(_01258_));
 sky130_fd_sc_hd__clkbuf_4 _10419_ (.A(_03388_),
    .X(_03422_));
 sky130_fd_sc_hd__mux2_1 _10420_ (.A0(\rbzero.tex_r1[17] ),
    .A1(\rbzero.tex_r1[18] ),
    .S(_03422_),
    .X(_03423_));
 sky130_fd_sc_hd__clkbuf_1 _10421_ (.A(_03423_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _10422_ (.A0(\rbzero.tex_r1[16] ),
    .A1(\rbzero.tex_r1[17] ),
    .S(_03422_),
    .X(_03424_));
 sky130_fd_sc_hd__clkbuf_1 _10423_ (.A(_03424_),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _10424_ (.A0(\rbzero.tex_r1[15] ),
    .A1(\rbzero.tex_r1[16] ),
    .S(_03422_),
    .X(_03425_));
 sky130_fd_sc_hd__clkbuf_1 _10425_ (.A(_03425_),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _10426_ (.A0(\rbzero.tex_r1[14] ),
    .A1(\rbzero.tex_r1[15] ),
    .S(_03422_),
    .X(_03426_));
 sky130_fd_sc_hd__clkbuf_1 _10427_ (.A(_03426_),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _10428_ (.A0(\rbzero.tex_r1[13] ),
    .A1(\rbzero.tex_r1[14] ),
    .S(_03422_),
    .X(_03427_));
 sky130_fd_sc_hd__clkbuf_1 _10429_ (.A(_03427_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _10430_ (.A0(\rbzero.tex_r1[12] ),
    .A1(\rbzero.tex_r1[13] ),
    .S(_03422_),
    .X(_03428_));
 sky130_fd_sc_hd__clkbuf_1 _10431_ (.A(_03428_),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _10432_ (.A0(\rbzero.tex_r1[11] ),
    .A1(\rbzero.tex_r1[12] ),
    .S(_03422_),
    .X(_03429_));
 sky130_fd_sc_hd__clkbuf_1 _10433_ (.A(_03429_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _10434_ (.A0(\rbzero.tex_r1[10] ),
    .A1(\rbzero.tex_r1[11] ),
    .S(_03422_),
    .X(_03430_));
 sky130_fd_sc_hd__clkbuf_1 _10435_ (.A(_03430_),
    .X(_01250_));
 sky130_fd_sc_hd__mux2_1 _10436_ (.A0(\rbzero.tex_r1[9] ),
    .A1(\rbzero.tex_r1[10] ),
    .S(_03422_),
    .X(_03431_));
 sky130_fd_sc_hd__clkbuf_1 _10437_ (.A(_03431_),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _10438_ (.A0(\rbzero.tex_r1[8] ),
    .A1(\rbzero.tex_r1[9] ),
    .S(_03422_),
    .X(_03432_));
 sky130_fd_sc_hd__clkbuf_1 _10439_ (.A(_03432_),
    .X(_01248_));
 sky130_fd_sc_hd__clkbuf_4 _10440_ (.A(_03388_),
    .X(_03433_));
 sky130_fd_sc_hd__mux2_1 _10441_ (.A0(\rbzero.tex_r1[7] ),
    .A1(\rbzero.tex_r1[8] ),
    .S(_03433_),
    .X(_03434_));
 sky130_fd_sc_hd__clkbuf_1 _10442_ (.A(_03434_),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _10443_ (.A0(\rbzero.tex_r1[6] ),
    .A1(\rbzero.tex_r1[7] ),
    .S(_03433_),
    .X(_03435_));
 sky130_fd_sc_hd__clkbuf_1 _10444_ (.A(_03435_),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _10445_ (.A0(\rbzero.tex_r1[5] ),
    .A1(\rbzero.tex_r1[6] ),
    .S(_03433_),
    .X(_03436_));
 sky130_fd_sc_hd__clkbuf_1 _10446_ (.A(_03436_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _10447_ (.A0(\rbzero.tex_r1[4] ),
    .A1(\rbzero.tex_r1[5] ),
    .S(_03433_),
    .X(_03437_));
 sky130_fd_sc_hd__clkbuf_1 _10448_ (.A(_03437_),
    .X(_01244_));
 sky130_fd_sc_hd__mux2_1 _10449_ (.A0(\rbzero.tex_r1[3] ),
    .A1(\rbzero.tex_r1[4] ),
    .S(_03433_),
    .X(_03438_));
 sky130_fd_sc_hd__clkbuf_1 _10450_ (.A(_03438_),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _10451_ (.A0(\rbzero.tex_r1[2] ),
    .A1(\rbzero.tex_r1[3] ),
    .S(_03433_),
    .X(_03439_));
 sky130_fd_sc_hd__clkbuf_1 _10452_ (.A(_03439_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _10453_ (.A0(\rbzero.tex_r1[1] ),
    .A1(\rbzero.tex_r1[2] ),
    .S(_03433_),
    .X(_03440_));
 sky130_fd_sc_hd__clkbuf_1 _10454_ (.A(_03440_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _10455_ (.A0(\rbzero.tex_r1[0] ),
    .A1(\rbzero.tex_r1[1] ),
    .S(_03433_),
    .X(_03441_));
 sky130_fd_sc_hd__clkbuf_1 _10456_ (.A(_03441_),
    .X(_01240_));
 sky130_fd_sc_hd__xnor2_4 _10457_ (.A(net46),
    .B(net45),
    .Y(_03442_));
 sky130_fd_sc_hd__nand2_1 _10458_ (.A(_03291_),
    .B(_03297_),
    .Y(_03443_));
 sky130_fd_sc_hd__or3_4 _10459_ (.A(_03289_),
    .B(_03442_),
    .C(_03443_),
    .X(_03444_));
 sky130_fd_sc_hd__clkbuf_4 _10460_ (.A(_03444_),
    .X(_03445_));
 sky130_fd_sc_hd__clkbuf_4 _10461_ (.A(_03445_),
    .X(_03446_));
 sky130_fd_sc_hd__mux2_1 _10462_ (.A0(net48),
    .A1(\rbzero.tex_r0[63] ),
    .S(_03446_),
    .X(_03447_));
 sky130_fd_sc_hd__clkbuf_1 _10463_ (.A(_03447_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _10464_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_03446_),
    .X(_03448_));
 sky130_fd_sc_hd__clkbuf_1 _10465_ (.A(_03448_),
    .X(_01238_));
 sky130_fd_sc_hd__mux2_1 _10466_ (.A0(\rbzero.tex_r0[62] ),
    .A1(\rbzero.tex_r0[61] ),
    .S(_03446_),
    .X(_03449_));
 sky130_fd_sc_hd__clkbuf_1 _10467_ (.A(_03449_),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _10468_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_03446_),
    .X(_03450_));
 sky130_fd_sc_hd__clkbuf_1 _10469_ (.A(_03450_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _10470_ (.A0(\rbzero.tex_r0[60] ),
    .A1(\rbzero.tex_r0[59] ),
    .S(_03446_),
    .X(_03451_));
 sky130_fd_sc_hd__clkbuf_1 _10471_ (.A(_03451_),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _10472_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(_03446_),
    .X(_03452_));
 sky130_fd_sc_hd__clkbuf_1 _10473_ (.A(_03452_),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _10474_ (.A0(\rbzero.tex_r0[58] ),
    .A1(\rbzero.tex_r0[57] ),
    .S(_03446_),
    .X(_03453_));
 sky130_fd_sc_hd__clkbuf_1 _10475_ (.A(_03453_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _10476_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(_03446_),
    .X(_03454_));
 sky130_fd_sc_hd__clkbuf_1 _10477_ (.A(_03454_),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _10478_ (.A0(\rbzero.tex_r0[56] ),
    .A1(\rbzero.tex_r0[55] ),
    .S(_03446_),
    .X(_03455_));
 sky130_fd_sc_hd__clkbuf_1 _10479_ (.A(_03455_),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _10480_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(_03446_),
    .X(_03456_));
 sky130_fd_sc_hd__clkbuf_1 _10481_ (.A(_03456_),
    .X(_01230_));
 sky130_fd_sc_hd__clkbuf_4 _10482_ (.A(_03445_),
    .X(_03457_));
 sky130_fd_sc_hd__mux2_1 _10483_ (.A0(\rbzero.tex_r0[54] ),
    .A1(\rbzero.tex_r0[53] ),
    .S(_03457_),
    .X(_03458_));
 sky130_fd_sc_hd__clkbuf_1 _10484_ (.A(_03458_),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _10485_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(_03457_),
    .X(_03459_));
 sky130_fd_sc_hd__clkbuf_1 _10486_ (.A(_03459_),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _10487_ (.A0(\rbzero.tex_r0[52] ),
    .A1(\rbzero.tex_r0[51] ),
    .S(_03457_),
    .X(_03460_));
 sky130_fd_sc_hd__clkbuf_1 _10488_ (.A(_03460_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _10489_ (.A0(\rbzero.tex_r0[51] ),
    .A1(\rbzero.tex_r0[50] ),
    .S(_03457_),
    .X(_03461_));
 sky130_fd_sc_hd__clkbuf_1 _10490_ (.A(_03461_),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _10491_ (.A0(\rbzero.tex_r0[50] ),
    .A1(\rbzero.tex_r0[49] ),
    .S(_03457_),
    .X(_03462_));
 sky130_fd_sc_hd__clkbuf_1 _10492_ (.A(_03462_),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _10493_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_03457_),
    .X(_03463_));
 sky130_fd_sc_hd__clkbuf_1 _10494_ (.A(_03463_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _10495_ (.A0(\rbzero.tex_r0[48] ),
    .A1(\rbzero.tex_r0[47] ),
    .S(_03457_),
    .X(_03464_));
 sky130_fd_sc_hd__clkbuf_1 _10496_ (.A(_03464_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _10497_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_03457_),
    .X(_03465_));
 sky130_fd_sc_hd__clkbuf_1 _10498_ (.A(_03465_),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _10499_ (.A0(\rbzero.tex_r0[46] ),
    .A1(\rbzero.tex_r0[45] ),
    .S(_03457_),
    .X(_03466_));
 sky130_fd_sc_hd__clkbuf_1 _10500_ (.A(_03466_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _10501_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_03457_),
    .X(_03467_));
 sky130_fd_sc_hd__clkbuf_1 _10502_ (.A(_03467_),
    .X(_01220_));
 sky130_fd_sc_hd__clkbuf_4 _10503_ (.A(_03445_),
    .X(_03468_));
 sky130_fd_sc_hd__mux2_1 _10504_ (.A0(\rbzero.tex_r0[44] ),
    .A1(\rbzero.tex_r0[43] ),
    .S(_03468_),
    .X(_03469_));
 sky130_fd_sc_hd__clkbuf_1 _10505_ (.A(_03469_),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _10506_ (.A0(\rbzero.tex_r0[43] ),
    .A1(\rbzero.tex_r0[42] ),
    .S(_03468_),
    .X(_03470_));
 sky130_fd_sc_hd__clkbuf_1 _10507_ (.A(_03470_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _10508_ (.A0(\rbzero.tex_r0[42] ),
    .A1(\rbzero.tex_r0[41] ),
    .S(_03468_),
    .X(_03471_));
 sky130_fd_sc_hd__clkbuf_1 _10509_ (.A(_03471_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _10510_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(_03468_),
    .X(_03472_));
 sky130_fd_sc_hd__clkbuf_1 _10511_ (.A(_03472_),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _10512_ (.A0(\rbzero.tex_r0[40] ),
    .A1(\rbzero.tex_r0[39] ),
    .S(_03468_),
    .X(_03473_));
 sky130_fd_sc_hd__clkbuf_1 _10513_ (.A(_03473_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _10514_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_03468_),
    .X(_03474_));
 sky130_fd_sc_hd__clkbuf_1 _10515_ (.A(_03474_),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _10516_ (.A0(\rbzero.tex_r0[38] ),
    .A1(\rbzero.tex_r0[37] ),
    .S(_03468_),
    .X(_03475_));
 sky130_fd_sc_hd__clkbuf_1 _10517_ (.A(_03475_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _10518_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_03468_),
    .X(_03476_));
 sky130_fd_sc_hd__clkbuf_1 _10519_ (.A(_03476_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _10520_ (.A0(\rbzero.tex_r0[36] ),
    .A1(\rbzero.tex_r0[35] ),
    .S(_03468_),
    .X(_03477_));
 sky130_fd_sc_hd__clkbuf_1 _10521_ (.A(_03477_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _10522_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(_03468_),
    .X(_03478_));
 sky130_fd_sc_hd__clkbuf_1 _10523_ (.A(_03478_),
    .X(_01210_));
 sky130_fd_sc_hd__clkbuf_4 _10524_ (.A(_03445_),
    .X(_03479_));
 sky130_fd_sc_hd__mux2_1 _10525_ (.A0(\rbzero.tex_r0[34] ),
    .A1(\rbzero.tex_r0[33] ),
    .S(_03479_),
    .X(_03480_));
 sky130_fd_sc_hd__clkbuf_1 _10526_ (.A(_03480_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _10527_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_03479_),
    .X(_03481_));
 sky130_fd_sc_hd__clkbuf_1 _10528_ (.A(_03481_),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _10529_ (.A0(\rbzero.tex_r0[32] ),
    .A1(\rbzero.tex_r0[31] ),
    .S(_03479_),
    .X(_03482_));
 sky130_fd_sc_hd__clkbuf_1 _10530_ (.A(_03482_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _10531_ (.A0(\rbzero.tex_r0[31] ),
    .A1(\rbzero.tex_r0[30] ),
    .S(_03479_),
    .X(_03483_));
 sky130_fd_sc_hd__clkbuf_1 _10532_ (.A(_03483_),
    .X(_01206_));
 sky130_fd_sc_hd__mux2_1 _10533_ (.A0(\rbzero.tex_r0[30] ),
    .A1(\rbzero.tex_r0[29] ),
    .S(_03479_),
    .X(_03484_));
 sky130_fd_sc_hd__clkbuf_1 _10534_ (.A(_03484_),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _10535_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_03479_),
    .X(_03485_));
 sky130_fd_sc_hd__clkbuf_1 _10536_ (.A(_03485_),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _10537_ (.A0(\rbzero.tex_r0[28] ),
    .A1(\rbzero.tex_r0[27] ),
    .S(_03479_),
    .X(_03486_));
 sky130_fd_sc_hd__clkbuf_1 _10538_ (.A(_03486_),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _10539_ (.A0(\rbzero.tex_r0[27] ),
    .A1(\rbzero.tex_r0[26] ),
    .S(_03479_),
    .X(_03487_));
 sky130_fd_sc_hd__clkbuf_1 _10540_ (.A(_03487_),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _10541_ (.A0(\rbzero.tex_r0[26] ),
    .A1(\rbzero.tex_r0[25] ),
    .S(_03479_),
    .X(_03488_));
 sky130_fd_sc_hd__clkbuf_1 _10542_ (.A(_03488_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _10543_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_03479_),
    .X(_03489_));
 sky130_fd_sc_hd__clkbuf_1 _10544_ (.A(_03489_),
    .X(_01200_));
 sky130_fd_sc_hd__clkbuf_4 _10545_ (.A(_03445_),
    .X(_03490_));
 sky130_fd_sc_hd__mux2_1 _10546_ (.A0(\rbzero.tex_r0[24] ),
    .A1(\rbzero.tex_r0[23] ),
    .S(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__clkbuf_1 _10547_ (.A(_03491_),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _10548_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(_03490_),
    .X(_03492_));
 sky130_fd_sc_hd__clkbuf_1 _10549_ (.A(_03492_),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _10550_ (.A0(\rbzero.tex_r0[22] ),
    .A1(\rbzero.tex_r0[21] ),
    .S(_03490_),
    .X(_03493_));
 sky130_fd_sc_hd__clkbuf_1 _10551_ (.A(_03493_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _10552_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(_03490_),
    .X(_03494_));
 sky130_fd_sc_hd__clkbuf_1 _10553_ (.A(_03494_),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _10554_ (.A0(\rbzero.tex_r0[20] ),
    .A1(\rbzero.tex_r0[19] ),
    .S(_03490_),
    .X(_03495_));
 sky130_fd_sc_hd__clkbuf_1 _10555_ (.A(_03495_),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _10556_ (.A0(\rbzero.tex_r0[19] ),
    .A1(\rbzero.tex_r0[18] ),
    .S(_03490_),
    .X(_03496_));
 sky130_fd_sc_hd__clkbuf_1 _10557_ (.A(_03496_),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _10558_ (.A0(\rbzero.tex_r0[18] ),
    .A1(\rbzero.tex_r0[17] ),
    .S(_03490_),
    .X(_03497_));
 sky130_fd_sc_hd__clkbuf_1 _10559_ (.A(_03497_),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _10560_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_03490_),
    .X(_03498_));
 sky130_fd_sc_hd__clkbuf_1 _10561_ (.A(_03498_),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _10562_ (.A0(\rbzero.tex_r0[16] ),
    .A1(\rbzero.tex_r0[15] ),
    .S(_03490_),
    .X(_03499_));
 sky130_fd_sc_hd__clkbuf_1 _10563_ (.A(_03499_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _10564_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(_03490_),
    .X(_03500_));
 sky130_fd_sc_hd__clkbuf_1 _10565_ (.A(_03500_),
    .X(_01190_));
 sky130_fd_sc_hd__clkbuf_4 _10566_ (.A(_03445_),
    .X(_03501_));
 sky130_fd_sc_hd__mux2_1 _10567_ (.A0(\rbzero.tex_r0[14] ),
    .A1(\rbzero.tex_r0[13] ),
    .S(_03501_),
    .X(_03502_));
 sky130_fd_sc_hd__clkbuf_1 _10568_ (.A(_03502_),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _10569_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(_03501_),
    .X(_03503_));
 sky130_fd_sc_hd__clkbuf_1 _10570_ (.A(_03503_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _10571_ (.A0(\rbzero.tex_r0[12] ),
    .A1(\rbzero.tex_r0[11] ),
    .S(_03501_),
    .X(_03504_));
 sky130_fd_sc_hd__clkbuf_1 _10572_ (.A(_03504_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _10573_ (.A0(\rbzero.tex_r0[11] ),
    .A1(\rbzero.tex_r0[10] ),
    .S(_03501_),
    .X(_03505_));
 sky130_fd_sc_hd__clkbuf_1 _10574_ (.A(_03505_),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _10575_ (.A0(\rbzero.tex_r0[10] ),
    .A1(\rbzero.tex_r0[9] ),
    .S(_03501_),
    .X(_03506_));
 sky130_fd_sc_hd__clkbuf_1 _10576_ (.A(_03506_),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _10577_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_03501_),
    .X(_03507_));
 sky130_fd_sc_hd__clkbuf_1 _10578_ (.A(_03507_),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _10579_ (.A0(\rbzero.tex_r0[8] ),
    .A1(\rbzero.tex_r0[7] ),
    .S(_03501_),
    .X(_03508_));
 sky130_fd_sc_hd__clkbuf_1 _10580_ (.A(_03508_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _10581_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_03501_),
    .X(_03509_));
 sky130_fd_sc_hd__clkbuf_1 _10582_ (.A(_03509_),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _10583_ (.A0(\rbzero.tex_r0[6] ),
    .A1(\rbzero.tex_r0[5] ),
    .S(_03501_),
    .X(_03510_));
 sky130_fd_sc_hd__clkbuf_1 _10584_ (.A(_03510_),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _10585_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_03501_),
    .X(_03511_));
 sky130_fd_sc_hd__clkbuf_1 _10586_ (.A(_03511_),
    .X(_01180_));
 sky130_fd_sc_hd__clkbuf_4 _10587_ (.A(_03445_),
    .X(_03512_));
 sky130_fd_sc_hd__mux2_1 _10588_ (.A0(\rbzero.tex_r0[4] ),
    .A1(\rbzero.tex_r0[3] ),
    .S(_03512_),
    .X(_03513_));
 sky130_fd_sc_hd__clkbuf_1 _10589_ (.A(_03513_),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _10590_ (.A0(\rbzero.tex_r0[3] ),
    .A1(\rbzero.tex_r0[2] ),
    .S(_03512_),
    .X(_03514_));
 sky130_fd_sc_hd__clkbuf_1 _10591_ (.A(_03514_),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _10592_ (.A0(\rbzero.tex_r0[2] ),
    .A1(\rbzero.tex_r0[1] ),
    .S(_03512_),
    .X(_03515_));
 sky130_fd_sc_hd__clkbuf_1 _10593_ (.A(_03515_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _10594_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_03512_),
    .X(_03516_));
 sky130_fd_sc_hd__clkbuf_1 _10595_ (.A(_03516_),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _10596_ (.A0(\rbzero.tex_g1[63] ),
    .A1(net49),
    .S(_03433_),
    .X(_03517_));
 sky130_fd_sc_hd__clkbuf_1 _10597_ (.A(_03517_),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _10598_ (.A0(\rbzero.tex_g1[62] ),
    .A1(\rbzero.tex_g1[63] ),
    .S(_03433_),
    .X(_03518_));
 sky130_fd_sc_hd__clkbuf_1 _10599_ (.A(_03518_),
    .X(_01174_));
 sky130_fd_sc_hd__clkbuf_4 _10600_ (.A(_03388_),
    .X(_03519_));
 sky130_fd_sc_hd__mux2_1 _10601_ (.A0(\rbzero.tex_g1[61] ),
    .A1(\rbzero.tex_g1[62] ),
    .S(_03519_),
    .X(_03520_));
 sky130_fd_sc_hd__clkbuf_1 _10602_ (.A(_03520_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _10603_ (.A0(\rbzero.tex_g1[60] ),
    .A1(\rbzero.tex_g1[61] ),
    .S(_03519_),
    .X(_03521_));
 sky130_fd_sc_hd__clkbuf_1 _10604_ (.A(_03521_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _10605_ (.A0(\rbzero.tex_g1[59] ),
    .A1(\rbzero.tex_g1[60] ),
    .S(_03519_),
    .X(_03522_));
 sky130_fd_sc_hd__clkbuf_1 _10606_ (.A(_03522_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _10607_ (.A0(\rbzero.tex_g1[58] ),
    .A1(\rbzero.tex_g1[59] ),
    .S(_03519_),
    .X(_03523_));
 sky130_fd_sc_hd__clkbuf_1 _10608_ (.A(_03523_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _10609_ (.A0(\rbzero.tex_g1[57] ),
    .A1(\rbzero.tex_g1[58] ),
    .S(_03519_),
    .X(_03524_));
 sky130_fd_sc_hd__clkbuf_1 _10610_ (.A(_03524_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _10611_ (.A0(\rbzero.tex_g1[56] ),
    .A1(\rbzero.tex_g1[57] ),
    .S(_03519_),
    .X(_03525_));
 sky130_fd_sc_hd__clkbuf_1 _10612_ (.A(_03525_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _10613_ (.A0(\rbzero.tex_g1[55] ),
    .A1(\rbzero.tex_g1[56] ),
    .S(_03519_),
    .X(_03526_));
 sky130_fd_sc_hd__clkbuf_1 _10614_ (.A(_03526_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _10615_ (.A0(\rbzero.tex_g1[54] ),
    .A1(\rbzero.tex_g1[55] ),
    .S(_03519_),
    .X(_03527_));
 sky130_fd_sc_hd__clkbuf_1 _10616_ (.A(_03527_),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _10617_ (.A0(\rbzero.tex_g1[53] ),
    .A1(\rbzero.tex_g1[54] ),
    .S(_03519_),
    .X(_03528_));
 sky130_fd_sc_hd__clkbuf_1 _10618_ (.A(_03528_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _10619_ (.A0(\rbzero.tex_g1[52] ),
    .A1(\rbzero.tex_g1[53] ),
    .S(_03519_),
    .X(_03529_));
 sky130_fd_sc_hd__clkbuf_1 _10620_ (.A(_03529_),
    .X(_01164_));
 sky130_fd_sc_hd__clkbuf_4 _10621_ (.A(_03388_),
    .X(_03530_));
 sky130_fd_sc_hd__mux2_1 _10622_ (.A0(\rbzero.tex_g1[51] ),
    .A1(\rbzero.tex_g1[52] ),
    .S(_03530_),
    .X(_03531_));
 sky130_fd_sc_hd__clkbuf_1 _10623_ (.A(_03531_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _10624_ (.A0(\rbzero.tex_g1[50] ),
    .A1(\rbzero.tex_g1[51] ),
    .S(_03530_),
    .X(_03532_));
 sky130_fd_sc_hd__clkbuf_1 _10625_ (.A(_03532_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _10626_ (.A0(\rbzero.tex_g1[49] ),
    .A1(\rbzero.tex_g1[50] ),
    .S(_03530_),
    .X(_03533_));
 sky130_fd_sc_hd__clkbuf_1 _10627_ (.A(_03533_),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(\rbzero.tex_g1[48] ),
    .A1(\rbzero.tex_g1[49] ),
    .S(_03530_),
    .X(_03534_));
 sky130_fd_sc_hd__clkbuf_1 _10629_ (.A(_03534_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _10630_ (.A0(\rbzero.tex_g1[47] ),
    .A1(\rbzero.tex_g1[48] ),
    .S(_03530_),
    .X(_03535_));
 sky130_fd_sc_hd__clkbuf_1 _10631_ (.A(_03535_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _10632_ (.A0(\rbzero.tex_g1[46] ),
    .A1(\rbzero.tex_g1[47] ),
    .S(_03530_),
    .X(_03536_));
 sky130_fd_sc_hd__clkbuf_1 _10633_ (.A(_03536_),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _10634_ (.A0(\rbzero.tex_g1[45] ),
    .A1(\rbzero.tex_g1[46] ),
    .S(_03530_),
    .X(_03537_));
 sky130_fd_sc_hd__clkbuf_1 _10635_ (.A(_03537_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _10636_ (.A0(\rbzero.tex_g1[44] ),
    .A1(\rbzero.tex_g1[45] ),
    .S(_03530_),
    .X(_03538_));
 sky130_fd_sc_hd__clkbuf_1 _10637_ (.A(_03538_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _10638_ (.A0(\rbzero.tex_g1[43] ),
    .A1(\rbzero.tex_g1[44] ),
    .S(_03530_),
    .X(_03539_));
 sky130_fd_sc_hd__clkbuf_1 _10639_ (.A(_03539_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _10640_ (.A0(\rbzero.tex_g1[42] ),
    .A1(\rbzero.tex_g1[43] ),
    .S(_03530_),
    .X(_03540_));
 sky130_fd_sc_hd__clkbuf_1 _10641_ (.A(_03540_),
    .X(_01154_));
 sky130_fd_sc_hd__clkbuf_4 _10642_ (.A(_03388_),
    .X(_03541_));
 sky130_fd_sc_hd__mux2_1 _10643_ (.A0(\rbzero.tex_g1[41] ),
    .A1(\rbzero.tex_g1[42] ),
    .S(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__clkbuf_1 _10644_ (.A(_03542_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(\rbzero.tex_g1[40] ),
    .A1(\rbzero.tex_g1[41] ),
    .S(_03541_),
    .X(_03543_));
 sky130_fd_sc_hd__clkbuf_1 _10646_ (.A(_03543_),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _10647_ (.A0(\rbzero.tex_g1[39] ),
    .A1(\rbzero.tex_g1[40] ),
    .S(_03541_),
    .X(_03544_));
 sky130_fd_sc_hd__clkbuf_1 _10648_ (.A(_03544_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _10649_ (.A0(\rbzero.tex_g1[38] ),
    .A1(\rbzero.tex_g1[39] ),
    .S(_03541_),
    .X(_03545_));
 sky130_fd_sc_hd__clkbuf_1 _10650_ (.A(_03545_),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _10651_ (.A0(\rbzero.tex_g1[37] ),
    .A1(\rbzero.tex_g1[38] ),
    .S(_03541_),
    .X(_03546_));
 sky130_fd_sc_hd__clkbuf_1 _10652_ (.A(_03546_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _10653_ (.A0(\rbzero.tex_g1[36] ),
    .A1(\rbzero.tex_g1[37] ),
    .S(_03541_),
    .X(_03547_));
 sky130_fd_sc_hd__clkbuf_1 _10654_ (.A(_03547_),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _10655_ (.A0(\rbzero.tex_g1[35] ),
    .A1(\rbzero.tex_g1[36] ),
    .S(_03541_),
    .X(_03548_));
 sky130_fd_sc_hd__clkbuf_1 _10656_ (.A(_03548_),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _10657_ (.A0(\rbzero.tex_g1[34] ),
    .A1(\rbzero.tex_g1[35] ),
    .S(_03541_),
    .X(_03549_));
 sky130_fd_sc_hd__clkbuf_1 _10658_ (.A(_03549_),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _10659_ (.A0(\rbzero.tex_g1[33] ),
    .A1(\rbzero.tex_g1[34] ),
    .S(_03541_),
    .X(_03550_));
 sky130_fd_sc_hd__clkbuf_1 _10660_ (.A(_03550_),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _10661_ (.A0(\rbzero.tex_g1[32] ),
    .A1(\rbzero.tex_g1[33] ),
    .S(_03541_),
    .X(_03551_));
 sky130_fd_sc_hd__clkbuf_1 _10662_ (.A(_03551_),
    .X(_01144_));
 sky130_fd_sc_hd__clkbuf_4 _10663_ (.A(_03388_),
    .X(_03552_));
 sky130_fd_sc_hd__mux2_1 _10664_ (.A0(\rbzero.tex_g1[31] ),
    .A1(\rbzero.tex_g1[32] ),
    .S(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__clkbuf_1 _10665_ (.A(_03553_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _10666_ (.A0(\rbzero.tex_g1[30] ),
    .A1(\rbzero.tex_g1[31] ),
    .S(_03552_),
    .X(_03554_));
 sky130_fd_sc_hd__clkbuf_1 _10667_ (.A(_03554_),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _10668_ (.A0(\rbzero.tex_g1[29] ),
    .A1(\rbzero.tex_g1[30] ),
    .S(_03552_),
    .X(_03555_));
 sky130_fd_sc_hd__clkbuf_1 _10669_ (.A(_03555_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _10670_ (.A0(\rbzero.tex_g1[28] ),
    .A1(\rbzero.tex_g1[29] ),
    .S(_03552_),
    .X(_03556_));
 sky130_fd_sc_hd__clkbuf_1 _10671_ (.A(_03556_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _10672_ (.A0(\rbzero.tex_g1[27] ),
    .A1(\rbzero.tex_g1[28] ),
    .S(_03552_),
    .X(_03557_));
 sky130_fd_sc_hd__clkbuf_1 _10673_ (.A(_03557_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _10674_ (.A0(\rbzero.tex_g1[26] ),
    .A1(\rbzero.tex_g1[27] ),
    .S(_03552_),
    .X(_03558_));
 sky130_fd_sc_hd__clkbuf_1 _10675_ (.A(_03558_),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _10676_ (.A0(\rbzero.tex_g1[25] ),
    .A1(\rbzero.tex_g1[26] ),
    .S(_03552_),
    .X(_03559_));
 sky130_fd_sc_hd__clkbuf_1 _10677_ (.A(_03559_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _10678_ (.A0(\rbzero.tex_g1[24] ),
    .A1(\rbzero.tex_g1[25] ),
    .S(_03552_),
    .X(_03560_));
 sky130_fd_sc_hd__clkbuf_1 _10679_ (.A(_03560_),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _10680_ (.A0(\rbzero.tex_g1[23] ),
    .A1(\rbzero.tex_g1[24] ),
    .S(_03552_),
    .X(_03561_));
 sky130_fd_sc_hd__clkbuf_1 _10681_ (.A(_03561_),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _10682_ (.A0(\rbzero.tex_g1[22] ),
    .A1(\rbzero.tex_g1[23] ),
    .S(_03552_),
    .X(_03562_));
 sky130_fd_sc_hd__clkbuf_1 _10683_ (.A(_03562_),
    .X(_01134_));
 sky130_fd_sc_hd__clkbuf_4 _10684_ (.A(_03388_),
    .X(_03563_));
 sky130_fd_sc_hd__mux2_1 _10685_ (.A0(\rbzero.tex_g1[21] ),
    .A1(\rbzero.tex_g1[22] ),
    .S(_03563_),
    .X(_03564_));
 sky130_fd_sc_hd__clkbuf_1 _10686_ (.A(_03564_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _10687_ (.A0(\rbzero.tex_g1[20] ),
    .A1(\rbzero.tex_g1[21] ),
    .S(_03563_),
    .X(_03565_));
 sky130_fd_sc_hd__clkbuf_1 _10688_ (.A(_03565_),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _10689_ (.A0(\rbzero.tex_g1[19] ),
    .A1(\rbzero.tex_g1[20] ),
    .S(_03563_),
    .X(_03566_));
 sky130_fd_sc_hd__clkbuf_1 _10690_ (.A(_03566_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _10691_ (.A0(\rbzero.tex_g1[18] ),
    .A1(\rbzero.tex_g1[19] ),
    .S(_03563_),
    .X(_03567_));
 sky130_fd_sc_hd__clkbuf_1 _10692_ (.A(_03567_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _10693_ (.A0(\rbzero.tex_g1[17] ),
    .A1(\rbzero.tex_g1[18] ),
    .S(_03563_),
    .X(_03568_));
 sky130_fd_sc_hd__clkbuf_1 _10694_ (.A(_03568_),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _10695_ (.A0(\rbzero.tex_g1[16] ),
    .A1(\rbzero.tex_g1[17] ),
    .S(_03563_),
    .X(_03569_));
 sky130_fd_sc_hd__clkbuf_1 _10696_ (.A(_03569_),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _10697_ (.A0(\rbzero.tex_g1[15] ),
    .A1(\rbzero.tex_g1[16] ),
    .S(_03563_),
    .X(_03570_));
 sky130_fd_sc_hd__clkbuf_1 _10698_ (.A(_03570_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _10699_ (.A0(\rbzero.tex_g1[14] ),
    .A1(\rbzero.tex_g1[15] ),
    .S(_03563_),
    .X(_03571_));
 sky130_fd_sc_hd__clkbuf_1 _10700_ (.A(_03571_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _10701_ (.A0(\rbzero.tex_g1[13] ),
    .A1(\rbzero.tex_g1[14] ),
    .S(_03563_),
    .X(_03572_));
 sky130_fd_sc_hd__clkbuf_1 _10702_ (.A(_03572_),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _10703_ (.A0(\rbzero.tex_g1[12] ),
    .A1(\rbzero.tex_g1[13] ),
    .S(_03563_),
    .X(_03573_));
 sky130_fd_sc_hd__clkbuf_1 _10704_ (.A(_03573_),
    .X(_01124_));
 sky130_fd_sc_hd__clkbuf_4 _10705_ (.A(_03298_),
    .X(_03574_));
 sky130_fd_sc_hd__mux2_1 _10706_ (.A0(\rbzero.tex_g1[11] ),
    .A1(\rbzero.tex_g1[12] ),
    .S(_03574_),
    .X(_03575_));
 sky130_fd_sc_hd__clkbuf_1 _10707_ (.A(_03575_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _10708_ (.A0(\rbzero.tex_g1[10] ),
    .A1(\rbzero.tex_g1[11] ),
    .S(_03574_),
    .X(_03576_));
 sky130_fd_sc_hd__clkbuf_1 _10709_ (.A(_03576_),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _10710_ (.A0(\rbzero.tex_g1[9] ),
    .A1(\rbzero.tex_g1[10] ),
    .S(_03574_),
    .X(_03577_));
 sky130_fd_sc_hd__clkbuf_1 _10711_ (.A(_03577_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _10712_ (.A0(\rbzero.tex_g1[8] ),
    .A1(\rbzero.tex_g1[9] ),
    .S(_03574_),
    .X(_03578_));
 sky130_fd_sc_hd__clkbuf_1 _10713_ (.A(_03578_),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _10714_ (.A0(\rbzero.tex_g1[7] ),
    .A1(\rbzero.tex_g1[8] ),
    .S(_03574_),
    .X(_03579_));
 sky130_fd_sc_hd__clkbuf_1 _10715_ (.A(_03579_),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _10716_ (.A0(\rbzero.tex_g1[6] ),
    .A1(\rbzero.tex_g1[7] ),
    .S(_03574_),
    .X(_03580_));
 sky130_fd_sc_hd__clkbuf_1 _10717_ (.A(_03580_),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _10718_ (.A0(\rbzero.tex_g1[5] ),
    .A1(\rbzero.tex_g1[6] ),
    .S(_03574_),
    .X(_03581_));
 sky130_fd_sc_hd__clkbuf_1 _10719_ (.A(_03581_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _10720_ (.A0(\rbzero.tex_g1[4] ),
    .A1(\rbzero.tex_g1[5] ),
    .S(_03574_),
    .X(_03582_));
 sky130_fd_sc_hd__clkbuf_1 _10721_ (.A(_03582_),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _10722_ (.A0(\rbzero.tex_g1[3] ),
    .A1(\rbzero.tex_g1[4] ),
    .S(_03574_),
    .X(_03583_));
 sky130_fd_sc_hd__clkbuf_1 _10723_ (.A(_03583_),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _10724_ (.A0(\rbzero.tex_g1[2] ),
    .A1(\rbzero.tex_g1[3] ),
    .S(_03574_),
    .X(_03584_));
 sky130_fd_sc_hd__clkbuf_1 _10725_ (.A(_03584_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _10726_ (.A0(\rbzero.tex_g1[1] ),
    .A1(\rbzero.tex_g1[2] ),
    .S(_03299_),
    .X(_03585_));
 sky130_fd_sc_hd__clkbuf_1 _10727_ (.A(_03585_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _10728_ (.A0(\rbzero.tex_g1[0] ),
    .A1(\rbzero.tex_g1[1] ),
    .S(_03299_),
    .X(_03586_));
 sky130_fd_sc_hd__clkbuf_1 _10729_ (.A(_03586_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _10730_ (.A0(net49),
    .A1(\rbzero.tex_g0[63] ),
    .S(_03512_),
    .X(_03587_));
 sky130_fd_sc_hd__clkbuf_1 _10731_ (.A(_03587_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _10732_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(_03512_),
    .X(_03588_));
 sky130_fd_sc_hd__clkbuf_1 _10733_ (.A(_03588_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _10734_ (.A0(\rbzero.tex_g0[62] ),
    .A1(\rbzero.tex_g0[61] ),
    .S(_03512_),
    .X(_03589_));
 sky130_fd_sc_hd__clkbuf_1 _10735_ (.A(_03589_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _10736_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_03512_),
    .X(_03590_));
 sky130_fd_sc_hd__clkbuf_1 _10737_ (.A(_03590_),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_1 _10738_ (.A0(\rbzero.tex_g0[60] ),
    .A1(\rbzero.tex_g0[59] ),
    .S(_03512_),
    .X(_03591_));
 sky130_fd_sc_hd__clkbuf_1 _10739_ (.A(_03591_),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _10740_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_03512_),
    .X(_03592_));
 sky130_fd_sc_hd__clkbuf_1 _10741_ (.A(_03592_),
    .X(_01106_));
 sky130_fd_sc_hd__clkbuf_4 _10742_ (.A(_03445_),
    .X(_03593_));
 sky130_fd_sc_hd__mux2_1 _10743_ (.A0(\rbzero.tex_g0[58] ),
    .A1(\rbzero.tex_g0[57] ),
    .S(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__clkbuf_1 _10744_ (.A(_03594_),
    .X(_01105_));
 sky130_fd_sc_hd__mux2_1 _10745_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(_03593_),
    .X(_03595_));
 sky130_fd_sc_hd__clkbuf_1 _10746_ (.A(_03595_),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_1 _10747_ (.A0(\rbzero.tex_g0[56] ),
    .A1(\rbzero.tex_g0[55] ),
    .S(_03593_),
    .X(_03596_));
 sky130_fd_sc_hd__clkbuf_1 _10748_ (.A(_03596_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _10749_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(_03593_),
    .X(_03597_));
 sky130_fd_sc_hd__clkbuf_1 _10750_ (.A(_03597_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _10751_ (.A0(\rbzero.tex_g0[54] ),
    .A1(\rbzero.tex_g0[53] ),
    .S(_03593_),
    .X(_03598_));
 sky130_fd_sc_hd__clkbuf_1 _10752_ (.A(_03598_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _10753_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(_03593_),
    .X(_03599_));
 sky130_fd_sc_hd__clkbuf_1 _10754_ (.A(_03599_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _10755_ (.A0(\rbzero.tex_g0[52] ),
    .A1(\rbzero.tex_g0[51] ),
    .S(_03593_),
    .X(_03600_));
 sky130_fd_sc_hd__clkbuf_1 _10756_ (.A(_03600_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _10757_ (.A0(\rbzero.tex_g0[51] ),
    .A1(\rbzero.tex_g0[50] ),
    .S(_03593_),
    .X(_03601_));
 sky130_fd_sc_hd__clkbuf_1 _10758_ (.A(_03601_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _10759_ (.A0(\rbzero.tex_g0[50] ),
    .A1(\rbzero.tex_g0[49] ),
    .S(_03593_),
    .X(_03602_));
 sky130_fd_sc_hd__clkbuf_1 _10760_ (.A(_03602_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _10761_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_03593_),
    .X(_03603_));
 sky130_fd_sc_hd__clkbuf_1 _10762_ (.A(_03603_),
    .X(_01096_));
 sky130_fd_sc_hd__clkbuf_4 _10763_ (.A(_03444_),
    .X(_03604_));
 sky130_fd_sc_hd__clkbuf_4 _10764_ (.A(_03604_),
    .X(_03605_));
 sky130_fd_sc_hd__mux2_1 _10765_ (.A0(\rbzero.tex_g0[48] ),
    .A1(\rbzero.tex_g0[47] ),
    .S(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__clkbuf_1 _10766_ (.A(_03606_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _10767_ (.A0(\rbzero.tex_g0[47] ),
    .A1(\rbzero.tex_g0[46] ),
    .S(_03605_),
    .X(_03607_));
 sky130_fd_sc_hd__clkbuf_1 _10768_ (.A(_03607_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _10769_ (.A0(\rbzero.tex_g0[46] ),
    .A1(\rbzero.tex_g0[45] ),
    .S(_03605_),
    .X(_03608_));
 sky130_fd_sc_hd__clkbuf_1 _10770_ (.A(_03608_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _10771_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(_03605_),
    .X(_03609_));
 sky130_fd_sc_hd__clkbuf_1 _10772_ (.A(_03609_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _10773_ (.A0(\rbzero.tex_g0[44] ),
    .A1(\rbzero.tex_g0[43] ),
    .S(_03605_),
    .X(_03610_));
 sky130_fd_sc_hd__clkbuf_1 _10774_ (.A(_03610_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _10775_ (.A0(\rbzero.tex_g0[43] ),
    .A1(\rbzero.tex_g0[42] ),
    .S(_03605_),
    .X(_03611_));
 sky130_fd_sc_hd__clkbuf_1 _10776_ (.A(_03611_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _10777_ (.A0(\rbzero.tex_g0[42] ),
    .A1(\rbzero.tex_g0[41] ),
    .S(_03605_),
    .X(_03612_));
 sky130_fd_sc_hd__clkbuf_1 _10778_ (.A(_03612_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_03605_),
    .X(_03613_));
 sky130_fd_sc_hd__clkbuf_1 _10780_ (.A(_03613_),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _10781_ (.A0(\rbzero.tex_g0[40] ),
    .A1(\rbzero.tex_g0[39] ),
    .S(_03605_),
    .X(_03614_));
 sky130_fd_sc_hd__clkbuf_1 _10782_ (.A(_03614_),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _10783_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_03605_),
    .X(_03615_));
 sky130_fd_sc_hd__clkbuf_1 _10784_ (.A(_03615_),
    .X(_01086_));
 sky130_fd_sc_hd__clkbuf_4 _10785_ (.A(_03604_),
    .X(_03616_));
 sky130_fd_sc_hd__mux2_1 _10786_ (.A0(\rbzero.tex_g0[38] ),
    .A1(\rbzero.tex_g0[37] ),
    .S(_03616_),
    .X(_03617_));
 sky130_fd_sc_hd__clkbuf_1 _10787_ (.A(_03617_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _10788_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_03616_),
    .X(_03618_));
 sky130_fd_sc_hd__clkbuf_1 _10789_ (.A(_03618_),
    .X(_01084_));
 sky130_fd_sc_hd__mux2_1 _10790_ (.A0(\rbzero.tex_g0[36] ),
    .A1(\rbzero.tex_g0[35] ),
    .S(_03616_),
    .X(_03619_));
 sky130_fd_sc_hd__clkbuf_1 _10791_ (.A(_03619_),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _10792_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(_03616_),
    .X(_03620_));
 sky130_fd_sc_hd__clkbuf_1 _10793_ (.A(_03620_),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _10794_ (.A0(\rbzero.tex_g0[34] ),
    .A1(\rbzero.tex_g0[33] ),
    .S(_03616_),
    .X(_03621_));
 sky130_fd_sc_hd__clkbuf_1 _10795_ (.A(_03621_),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _10796_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_03616_),
    .X(_03622_));
 sky130_fd_sc_hd__clkbuf_1 _10797_ (.A(_03622_),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _10798_ (.A0(\rbzero.tex_g0[32] ),
    .A1(\rbzero.tex_g0[31] ),
    .S(_03616_),
    .X(_03623_));
 sky130_fd_sc_hd__clkbuf_1 _10799_ (.A(_03623_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _10800_ (.A0(\rbzero.tex_g0[31] ),
    .A1(\rbzero.tex_g0[30] ),
    .S(_03616_),
    .X(_03624_));
 sky130_fd_sc_hd__clkbuf_1 _10801_ (.A(_03624_),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _10802_ (.A0(\rbzero.tex_g0[30] ),
    .A1(\rbzero.tex_g0[29] ),
    .S(_03616_),
    .X(_03625_));
 sky130_fd_sc_hd__clkbuf_1 _10803_ (.A(_03625_),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _10804_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_03616_),
    .X(_03626_));
 sky130_fd_sc_hd__clkbuf_1 _10805_ (.A(_03626_),
    .X(_01076_));
 sky130_fd_sc_hd__clkbuf_4 _10806_ (.A(_03604_),
    .X(_03627_));
 sky130_fd_sc_hd__mux2_1 _10807_ (.A0(\rbzero.tex_g0[28] ),
    .A1(\rbzero.tex_g0[27] ),
    .S(_03627_),
    .X(_03628_));
 sky130_fd_sc_hd__clkbuf_1 _10808_ (.A(_03628_),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _10809_ (.A0(\rbzero.tex_g0[27] ),
    .A1(\rbzero.tex_g0[26] ),
    .S(_03627_),
    .X(_03629_));
 sky130_fd_sc_hd__clkbuf_1 _10810_ (.A(_03629_),
    .X(_01074_));
 sky130_fd_sc_hd__mux2_1 _10811_ (.A0(\rbzero.tex_g0[26] ),
    .A1(\rbzero.tex_g0[25] ),
    .S(_03627_),
    .X(_03630_));
 sky130_fd_sc_hd__clkbuf_1 _10812_ (.A(_03630_),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _10813_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_03627_),
    .X(_03631_));
 sky130_fd_sc_hd__clkbuf_1 _10814_ (.A(_03631_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _10815_ (.A0(\rbzero.tex_g0[24] ),
    .A1(\rbzero.tex_g0[23] ),
    .S(_03627_),
    .X(_03632_));
 sky130_fd_sc_hd__clkbuf_1 _10816_ (.A(_03632_),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _10817_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(_03627_),
    .X(_03633_));
 sky130_fd_sc_hd__clkbuf_1 _10818_ (.A(_03633_),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _10819_ (.A0(\rbzero.tex_g0[22] ),
    .A1(\rbzero.tex_g0[21] ),
    .S(_03627_),
    .X(_03634_));
 sky130_fd_sc_hd__clkbuf_1 _10820_ (.A(_03634_),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _10821_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(_03627_),
    .X(_03635_));
 sky130_fd_sc_hd__clkbuf_1 _10822_ (.A(_03635_),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _10823_ (.A0(\rbzero.tex_g0[20] ),
    .A1(\rbzero.tex_g0[19] ),
    .S(_03627_),
    .X(_03636_));
 sky130_fd_sc_hd__clkbuf_1 _10824_ (.A(_03636_),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _10825_ (.A0(\rbzero.tex_g0[19] ),
    .A1(\rbzero.tex_g0[18] ),
    .S(_03627_),
    .X(_03637_));
 sky130_fd_sc_hd__clkbuf_1 _10826_ (.A(_03637_),
    .X(_01066_));
 sky130_fd_sc_hd__clkbuf_4 _10827_ (.A(_03604_),
    .X(_03638_));
 sky130_fd_sc_hd__mux2_1 _10828_ (.A0(\rbzero.tex_g0[18] ),
    .A1(\rbzero.tex_g0[17] ),
    .S(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__clkbuf_1 _10829_ (.A(_03639_),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_1 _10830_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_03638_),
    .X(_03640_));
 sky130_fd_sc_hd__clkbuf_1 _10831_ (.A(_03640_),
    .X(_01064_));
 sky130_fd_sc_hd__mux2_1 _10832_ (.A0(\rbzero.tex_g0[16] ),
    .A1(\rbzero.tex_g0[15] ),
    .S(_03638_),
    .X(_03641_));
 sky130_fd_sc_hd__clkbuf_1 _10833_ (.A(_03641_),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _10834_ (.A0(\rbzero.tex_g0[15] ),
    .A1(\rbzero.tex_g0[14] ),
    .S(_03638_),
    .X(_03642_));
 sky130_fd_sc_hd__clkbuf_1 _10835_ (.A(_03642_),
    .X(_01062_));
 sky130_fd_sc_hd__mux2_1 _10836_ (.A0(\rbzero.tex_g0[14] ),
    .A1(\rbzero.tex_g0[13] ),
    .S(_03638_),
    .X(_03643_));
 sky130_fd_sc_hd__clkbuf_1 _10837_ (.A(_03643_),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _10838_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_03638_),
    .X(_03644_));
 sky130_fd_sc_hd__clkbuf_1 _10839_ (.A(_03644_),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_1 _10840_ (.A0(\rbzero.tex_g0[12] ),
    .A1(\rbzero.tex_g0[11] ),
    .S(_03638_),
    .X(_03645_));
 sky130_fd_sc_hd__clkbuf_1 _10841_ (.A(_03645_),
    .X(_01059_));
 sky130_fd_sc_hd__mux2_1 _10842_ (.A0(\rbzero.tex_g0[11] ),
    .A1(\rbzero.tex_g0[10] ),
    .S(_03638_),
    .X(_03646_));
 sky130_fd_sc_hd__clkbuf_1 _10843_ (.A(_03646_),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _10844_ (.A0(\rbzero.tex_g0[10] ),
    .A1(\rbzero.tex_g0[9] ),
    .S(_03638_),
    .X(_03647_));
 sky130_fd_sc_hd__clkbuf_1 _10845_ (.A(_03647_),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_1 _10846_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_03638_),
    .X(_03648_));
 sky130_fd_sc_hd__clkbuf_1 _10847_ (.A(_03648_),
    .X(_01056_));
 sky130_fd_sc_hd__clkbuf_4 _10848_ (.A(_03604_),
    .X(_03649_));
 sky130_fd_sc_hd__mux2_1 _10849_ (.A0(\rbzero.tex_g0[8] ),
    .A1(\rbzero.tex_g0[7] ),
    .S(_03649_),
    .X(_03650_));
 sky130_fd_sc_hd__clkbuf_1 _10850_ (.A(_03650_),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _10851_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(_03649_),
    .X(_03651_));
 sky130_fd_sc_hd__clkbuf_1 _10852_ (.A(_03651_),
    .X(_01054_));
 sky130_fd_sc_hd__mux2_1 _10853_ (.A0(\rbzero.tex_g0[6] ),
    .A1(\rbzero.tex_g0[5] ),
    .S(_03649_),
    .X(_03652_));
 sky130_fd_sc_hd__clkbuf_1 _10854_ (.A(_03652_),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _10855_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_03649_),
    .X(_03653_));
 sky130_fd_sc_hd__clkbuf_1 _10856_ (.A(_03653_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _10857_ (.A0(\rbzero.tex_g0[4] ),
    .A1(\rbzero.tex_g0[3] ),
    .S(_03649_),
    .X(_03654_));
 sky130_fd_sc_hd__clkbuf_1 _10858_ (.A(_03654_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _10859_ (.A0(\rbzero.tex_g0[3] ),
    .A1(\rbzero.tex_g0[2] ),
    .S(_03649_),
    .X(_03655_));
 sky130_fd_sc_hd__clkbuf_1 _10860_ (.A(_03655_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _10861_ (.A0(\rbzero.tex_g0[2] ),
    .A1(\rbzero.tex_g0[1] ),
    .S(_03649_),
    .X(_03656_));
 sky130_fd_sc_hd__clkbuf_1 _10862_ (.A(_03656_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _10863_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_03649_),
    .X(_03657_));
 sky130_fd_sc_hd__clkbuf_1 _10864_ (.A(_03657_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _10865_ (.A0(net50),
    .A1(\rbzero.tex_b0[63] ),
    .S(_03649_),
    .X(_03658_));
 sky130_fd_sc_hd__clkbuf_1 _10866_ (.A(_03658_),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _10867_ (.A0(\rbzero.tex_b0[63] ),
    .A1(\rbzero.tex_b0[62] ),
    .S(_03649_),
    .X(_03659_));
 sky130_fd_sc_hd__clkbuf_1 _10868_ (.A(_03659_),
    .X(_00877_));
 sky130_fd_sc_hd__clkbuf_4 _10869_ (.A(_03604_),
    .X(_03660_));
 sky130_fd_sc_hd__mux2_1 _10870_ (.A0(\rbzero.tex_b0[62] ),
    .A1(\rbzero.tex_b0[61] ),
    .S(_03660_),
    .X(_03661_));
 sky130_fd_sc_hd__clkbuf_1 _10871_ (.A(_03661_),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _10872_ (.A0(\rbzero.tex_b0[61] ),
    .A1(\rbzero.tex_b0[60] ),
    .S(_03660_),
    .X(_03662_));
 sky130_fd_sc_hd__clkbuf_1 _10873_ (.A(_03662_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _10874_ (.A0(\rbzero.tex_b0[60] ),
    .A1(\rbzero.tex_b0[59] ),
    .S(_03660_),
    .X(_03663_));
 sky130_fd_sc_hd__clkbuf_1 _10875_ (.A(_03663_),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _10876_ (.A0(\rbzero.tex_b0[59] ),
    .A1(\rbzero.tex_b0[58] ),
    .S(_03660_),
    .X(_03664_));
 sky130_fd_sc_hd__clkbuf_1 _10877_ (.A(_03664_),
    .X(_00873_));
 sky130_fd_sc_hd__mux2_1 _10878_ (.A0(\rbzero.tex_b0[58] ),
    .A1(\rbzero.tex_b0[57] ),
    .S(_03660_),
    .X(_03665_));
 sky130_fd_sc_hd__clkbuf_1 _10879_ (.A(_03665_),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _10880_ (.A0(\rbzero.tex_b0[57] ),
    .A1(\rbzero.tex_b0[56] ),
    .S(_03660_),
    .X(_03666_));
 sky130_fd_sc_hd__clkbuf_1 _10881_ (.A(_03666_),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _10882_ (.A0(\rbzero.tex_b0[56] ),
    .A1(\rbzero.tex_b0[55] ),
    .S(_03660_),
    .X(_03667_));
 sky130_fd_sc_hd__clkbuf_1 _10883_ (.A(_03667_),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _10884_ (.A0(\rbzero.tex_b0[55] ),
    .A1(\rbzero.tex_b0[54] ),
    .S(_03660_),
    .X(_03668_));
 sky130_fd_sc_hd__clkbuf_1 _10885_ (.A(_03668_),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _10886_ (.A0(\rbzero.tex_b0[54] ),
    .A1(\rbzero.tex_b0[53] ),
    .S(_03660_),
    .X(_03669_));
 sky130_fd_sc_hd__clkbuf_1 _10887_ (.A(_03669_),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _10888_ (.A0(\rbzero.tex_b0[53] ),
    .A1(\rbzero.tex_b0[52] ),
    .S(_03660_),
    .X(_03670_));
 sky130_fd_sc_hd__clkbuf_1 _10889_ (.A(_03670_),
    .X(_00867_));
 sky130_fd_sc_hd__clkbuf_4 _10890_ (.A(_03604_),
    .X(_03671_));
 sky130_fd_sc_hd__mux2_1 _10891_ (.A0(\rbzero.tex_b0[52] ),
    .A1(\rbzero.tex_b0[51] ),
    .S(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__clkbuf_1 _10892_ (.A(_03672_),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _10893_ (.A0(\rbzero.tex_b0[51] ),
    .A1(\rbzero.tex_b0[50] ),
    .S(_03671_),
    .X(_03673_));
 sky130_fd_sc_hd__clkbuf_1 _10894_ (.A(_03673_),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _10895_ (.A0(\rbzero.tex_b0[50] ),
    .A1(\rbzero.tex_b0[49] ),
    .S(_03671_),
    .X(_03674_));
 sky130_fd_sc_hd__clkbuf_1 _10896_ (.A(_03674_),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(\rbzero.tex_b0[49] ),
    .A1(\rbzero.tex_b0[48] ),
    .S(_03671_),
    .X(_03675_));
 sky130_fd_sc_hd__clkbuf_1 _10898_ (.A(_03675_),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _10899_ (.A0(\rbzero.tex_b0[48] ),
    .A1(\rbzero.tex_b0[47] ),
    .S(_03671_),
    .X(_03676_));
 sky130_fd_sc_hd__clkbuf_1 _10900_ (.A(_03676_),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_1 _10901_ (.A0(\rbzero.tex_b0[47] ),
    .A1(\rbzero.tex_b0[46] ),
    .S(_03671_),
    .X(_03677_));
 sky130_fd_sc_hd__clkbuf_1 _10902_ (.A(_03677_),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _10903_ (.A0(\rbzero.tex_b0[46] ),
    .A1(\rbzero.tex_b0[45] ),
    .S(_03671_),
    .X(_03678_));
 sky130_fd_sc_hd__clkbuf_1 _10904_ (.A(_03678_),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _10905_ (.A0(\rbzero.tex_b0[45] ),
    .A1(\rbzero.tex_b0[44] ),
    .S(_03671_),
    .X(_03679_));
 sky130_fd_sc_hd__clkbuf_1 _10906_ (.A(_03679_),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _10907_ (.A0(\rbzero.tex_b0[44] ),
    .A1(\rbzero.tex_b0[43] ),
    .S(_03671_),
    .X(_03680_));
 sky130_fd_sc_hd__clkbuf_1 _10908_ (.A(_03680_),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _10909_ (.A0(\rbzero.tex_b0[43] ),
    .A1(\rbzero.tex_b0[42] ),
    .S(_03671_),
    .X(_03681_));
 sky130_fd_sc_hd__clkbuf_1 _10910_ (.A(_03681_),
    .X(_00857_));
 sky130_fd_sc_hd__clkbuf_4 _10911_ (.A(_03604_),
    .X(_03682_));
 sky130_fd_sc_hd__mux2_1 _10912_ (.A0(\rbzero.tex_b0[42] ),
    .A1(\rbzero.tex_b0[41] ),
    .S(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__clkbuf_1 _10913_ (.A(_03683_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _10914_ (.A0(\rbzero.tex_b0[41] ),
    .A1(\rbzero.tex_b0[40] ),
    .S(_03682_),
    .X(_03684_));
 sky130_fd_sc_hd__clkbuf_1 _10915_ (.A(_03684_),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _10916_ (.A0(\rbzero.tex_b0[40] ),
    .A1(\rbzero.tex_b0[39] ),
    .S(_03682_),
    .X(_03685_));
 sky130_fd_sc_hd__clkbuf_1 _10917_ (.A(_03685_),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _10918_ (.A0(\rbzero.tex_b0[39] ),
    .A1(\rbzero.tex_b0[38] ),
    .S(_03682_),
    .X(_03686_));
 sky130_fd_sc_hd__clkbuf_1 _10919_ (.A(_03686_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _10920_ (.A0(\rbzero.tex_b0[38] ),
    .A1(\rbzero.tex_b0[37] ),
    .S(_03682_),
    .X(_03687_));
 sky130_fd_sc_hd__clkbuf_1 _10921_ (.A(_03687_),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _10922_ (.A0(\rbzero.tex_b0[37] ),
    .A1(\rbzero.tex_b0[36] ),
    .S(_03682_),
    .X(_03688_));
 sky130_fd_sc_hd__clkbuf_1 _10923_ (.A(_03688_),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _10924_ (.A0(\rbzero.tex_b0[36] ),
    .A1(\rbzero.tex_b0[35] ),
    .S(_03682_),
    .X(_03689_));
 sky130_fd_sc_hd__clkbuf_1 _10925_ (.A(_03689_),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _10926_ (.A0(\rbzero.tex_b0[35] ),
    .A1(\rbzero.tex_b0[34] ),
    .S(_03682_),
    .X(_03690_));
 sky130_fd_sc_hd__clkbuf_1 _10927_ (.A(_03690_),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _10928_ (.A0(\rbzero.tex_b0[34] ),
    .A1(\rbzero.tex_b0[33] ),
    .S(_03682_),
    .X(_03691_));
 sky130_fd_sc_hd__clkbuf_1 _10929_ (.A(_03691_),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _10930_ (.A0(\rbzero.tex_b0[33] ),
    .A1(\rbzero.tex_b0[32] ),
    .S(_03682_),
    .X(_03692_));
 sky130_fd_sc_hd__clkbuf_1 _10931_ (.A(_03692_),
    .X(_00847_));
 sky130_fd_sc_hd__clkbuf_4 _10932_ (.A(_03604_),
    .X(_03693_));
 sky130_fd_sc_hd__mux2_1 _10933_ (.A0(\rbzero.tex_b0[32] ),
    .A1(\rbzero.tex_b0[31] ),
    .S(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__clkbuf_1 _10934_ (.A(_03694_),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _10935_ (.A0(\rbzero.tex_b0[31] ),
    .A1(\rbzero.tex_b0[30] ),
    .S(_03693_),
    .X(_03695_));
 sky130_fd_sc_hd__clkbuf_1 _10936_ (.A(_03695_),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _10937_ (.A0(\rbzero.tex_b0[30] ),
    .A1(\rbzero.tex_b0[29] ),
    .S(_03693_),
    .X(_03696_));
 sky130_fd_sc_hd__clkbuf_1 _10938_ (.A(_03696_),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _10939_ (.A0(\rbzero.tex_b0[29] ),
    .A1(\rbzero.tex_b0[28] ),
    .S(_03693_),
    .X(_03697_));
 sky130_fd_sc_hd__clkbuf_1 _10940_ (.A(_03697_),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _10941_ (.A0(\rbzero.tex_b0[28] ),
    .A1(\rbzero.tex_b0[27] ),
    .S(_03693_),
    .X(_03698_));
 sky130_fd_sc_hd__clkbuf_1 _10942_ (.A(_03698_),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _10943_ (.A0(\rbzero.tex_b0[27] ),
    .A1(\rbzero.tex_b0[26] ),
    .S(_03693_),
    .X(_03699_));
 sky130_fd_sc_hd__clkbuf_1 _10944_ (.A(_03699_),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _10945_ (.A0(\rbzero.tex_b0[26] ),
    .A1(\rbzero.tex_b0[25] ),
    .S(_03693_),
    .X(_03700_));
 sky130_fd_sc_hd__clkbuf_1 _10946_ (.A(_03700_),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _10947_ (.A0(\rbzero.tex_b0[25] ),
    .A1(\rbzero.tex_b0[24] ),
    .S(_03693_),
    .X(_03701_));
 sky130_fd_sc_hd__clkbuf_1 _10948_ (.A(_03701_),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _10949_ (.A0(\rbzero.tex_b0[24] ),
    .A1(\rbzero.tex_b0[23] ),
    .S(_03693_),
    .X(_03702_));
 sky130_fd_sc_hd__clkbuf_1 _10950_ (.A(_03702_),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _10951_ (.A0(\rbzero.tex_b0[23] ),
    .A1(\rbzero.tex_b0[22] ),
    .S(_03693_),
    .X(_03703_));
 sky130_fd_sc_hd__clkbuf_1 _10952_ (.A(_03703_),
    .X(_00837_));
 sky130_fd_sc_hd__clkbuf_4 _10953_ (.A(_03604_),
    .X(_03704_));
 sky130_fd_sc_hd__mux2_1 _10954_ (.A0(\rbzero.tex_b0[22] ),
    .A1(\rbzero.tex_b0[21] ),
    .S(_03704_),
    .X(_03705_));
 sky130_fd_sc_hd__clkbuf_1 _10955_ (.A(_03705_),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _10956_ (.A0(\rbzero.tex_b0[21] ),
    .A1(\rbzero.tex_b0[20] ),
    .S(_03704_),
    .X(_03706_));
 sky130_fd_sc_hd__clkbuf_1 _10957_ (.A(_03706_),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _10958_ (.A0(\rbzero.tex_b0[20] ),
    .A1(\rbzero.tex_b0[19] ),
    .S(_03704_),
    .X(_03707_));
 sky130_fd_sc_hd__clkbuf_1 _10959_ (.A(_03707_),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _10960_ (.A0(\rbzero.tex_b0[19] ),
    .A1(\rbzero.tex_b0[18] ),
    .S(_03704_),
    .X(_03708_));
 sky130_fd_sc_hd__clkbuf_1 _10961_ (.A(_03708_),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_1 _10962_ (.A0(\rbzero.tex_b0[18] ),
    .A1(\rbzero.tex_b0[17] ),
    .S(_03704_),
    .X(_03709_));
 sky130_fd_sc_hd__clkbuf_1 _10963_ (.A(_03709_),
    .X(_00832_));
 sky130_fd_sc_hd__mux2_1 _10964_ (.A0(\rbzero.tex_b0[17] ),
    .A1(\rbzero.tex_b0[16] ),
    .S(_03704_),
    .X(_03710_));
 sky130_fd_sc_hd__clkbuf_1 _10965_ (.A(_03710_),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _10966_ (.A0(\rbzero.tex_b0[16] ),
    .A1(\rbzero.tex_b0[15] ),
    .S(_03704_),
    .X(_03711_));
 sky130_fd_sc_hd__clkbuf_1 _10967_ (.A(_03711_),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _10968_ (.A0(\rbzero.tex_b0[15] ),
    .A1(\rbzero.tex_b0[14] ),
    .S(_03704_),
    .X(_03712_));
 sky130_fd_sc_hd__clkbuf_1 _10969_ (.A(_03712_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _10970_ (.A0(\rbzero.tex_b0[14] ),
    .A1(\rbzero.tex_b0[13] ),
    .S(_03704_),
    .X(_03713_));
 sky130_fd_sc_hd__clkbuf_1 _10971_ (.A(_03713_),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _10972_ (.A0(\rbzero.tex_b0[13] ),
    .A1(\rbzero.tex_b0[12] ),
    .S(_03704_),
    .X(_03714_));
 sky130_fd_sc_hd__clkbuf_1 _10973_ (.A(_03714_),
    .X(_00827_));
 sky130_fd_sc_hd__clkbuf_4 _10974_ (.A(_03444_),
    .X(_03715_));
 sky130_fd_sc_hd__mux2_1 _10975_ (.A0(\rbzero.tex_b0[12] ),
    .A1(\rbzero.tex_b0[11] ),
    .S(_03715_),
    .X(_03716_));
 sky130_fd_sc_hd__clkbuf_1 _10976_ (.A(_03716_),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _10977_ (.A0(\rbzero.tex_b0[11] ),
    .A1(\rbzero.tex_b0[10] ),
    .S(_03715_),
    .X(_03717_));
 sky130_fd_sc_hd__clkbuf_1 _10978_ (.A(_03717_),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _10979_ (.A0(\rbzero.tex_b0[10] ),
    .A1(\rbzero.tex_b0[9] ),
    .S(_03715_),
    .X(_03718_));
 sky130_fd_sc_hd__clkbuf_1 _10980_ (.A(_03718_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _10981_ (.A0(\rbzero.tex_b0[9] ),
    .A1(\rbzero.tex_b0[8] ),
    .S(_03715_),
    .X(_03719_));
 sky130_fd_sc_hd__clkbuf_1 _10982_ (.A(_03719_),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _10983_ (.A0(\rbzero.tex_b0[8] ),
    .A1(\rbzero.tex_b0[7] ),
    .S(_03715_),
    .X(_03720_));
 sky130_fd_sc_hd__clkbuf_1 _10984_ (.A(_03720_),
    .X(_00822_));
 sky130_fd_sc_hd__mux2_1 _10985_ (.A0(\rbzero.tex_b0[7] ),
    .A1(\rbzero.tex_b0[6] ),
    .S(_03715_),
    .X(_03721_));
 sky130_fd_sc_hd__clkbuf_1 _10986_ (.A(_03721_),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _10987_ (.A0(\rbzero.tex_b0[6] ),
    .A1(\rbzero.tex_b0[5] ),
    .S(_03715_),
    .X(_03722_));
 sky130_fd_sc_hd__clkbuf_1 _10988_ (.A(_03722_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _10989_ (.A0(\rbzero.tex_b0[5] ),
    .A1(\rbzero.tex_b0[4] ),
    .S(_03715_),
    .X(_03723_));
 sky130_fd_sc_hd__clkbuf_1 _10990_ (.A(_03723_),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_1 _10991_ (.A0(\rbzero.tex_b0[4] ),
    .A1(\rbzero.tex_b0[3] ),
    .S(_03715_),
    .X(_03724_));
 sky130_fd_sc_hd__clkbuf_1 _10992_ (.A(_03724_),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_1 _10993_ (.A0(\rbzero.tex_b0[3] ),
    .A1(\rbzero.tex_b0[2] ),
    .S(_03715_),
    .X(_03725_));
 sky130_fd_sc_hd__clkbuf_1 _10994_ (.A(_03725_),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_1 _10995_ (.A0(\rbzero.tex_b0[2] ),
    .A1(\rbzero.tex_b0[1] ),
    .S(_03445_),
    .X(_03726_));
 sky130_fd_sc_hd__clkbuf_1 _10996_ (.A(_03726_),
    .X(_00816_));
 sky130_fd_sc_hd__mux2_1 _10997_ (.A0(\rbzero.tex_b0[1] ),
    .A1(\rbzero.tex_b0[0] ),
    .S(_03445_),
    .X(_03727_));
 sky130_fd_sc_hd__clkbuf_1 _10998_ (.A(_03727_),
    .X(_00815_));
 sky130_fd_sc_hd__clkinv_4 _10999_ (.A(\rbzero.vga_sync.vsync ),
    .Y(o_vsync));
 sky130_fd_sc_hd__nand2_1 _11000_ (.A(o_vsync),
    .B(_03292_),
    .Y(_03728_));
 sky130_fd_sc_hd__buf_4 _11001_ (.A(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__buf_4 _11002_ (.A(_03729_),
    .X(_03730_));
 sky130_fd_sc_hd__inv_2 _11003_ (.A(\rbzero.wall_tracer.state[1] ),
    .Y(_03731_));
 sky130_fd_sc_hd__inv_2 _11004_ (.A(\rbzero.map_rom.i_row[4] ),
    .Y(_03732_));
 sky130_fd_sc_hd__buf_2 _11005_ (.A(\rbzero.map_rom.b6 ),
    .X(_03733_));
 sky130_fd_sc_hd__nand2_1 _11006_ (.A(_03733_),
    .B(\rbzero.map_rom.a6 ),
    .Y(_03734_));
 sky130_fd_sc_hd__inv_2 _11007_ (.A(\rbzero.map_rom.f3 ),
    .Y(_03735_));
 sky130_fd_sc_hd__clkbuf_4 _11008_ (.A(\rbzero.map_rom.f2 ),
    .X(_03736_));
 sky130_fd_sc_hd__inv_2 _11009_ (.A(_03736_),
    .Y(_03737_));
 sky130_fd_sc_hd__or3b_1 _11010_ (.A(_03735_),
    .B(_03737_),
    .C_N(_03733_),
    .X(_03738_));
 sky130_fd_sc_hd__o21ai_1 _11011_ (.A1(_03732_),
    .A2(_03734_),
    .B1(_03738_),
    .Y(_03739_));
 sky130_fd_sc_hd__xor2_1 _11012_ (.A(_03736_),
    .B(_03733_),
    .X(_03740_));
 sky130_fd_sc_hd__nand2_1 _11013_ (.A(\rbzero.map_rom.f3 ),
    .B(\rbzero.map_rom.c6 ),
    .Y(_03741_));
 sky130_fd_sc_hd__inv_2 _11014_ (.A(\rbzero.map_rom.f4 ),
    .Y(_03742_));
 sky130_fd_sc_hd__inv_2 _11015_ (.A(\rbzero.map_rom.d6 ),
    .Y(_03743_));
 sky130_fd_sc_hd__inv_2 _11016_ (.A(\rbzero.map_rom.a6 ),
    .Y(_03744_));
 sky130_fd_sc_hd__o22a_1 _11017_ (.A1(\rbzero.map_rom.f4 ),
    .A2(\rbzero.map_rom.d6 ),
    .B1(\rbzero.map_rom.c6 ),
    .B2(\rbzero.map_rom.f3 ),
    .X(_03745_));
 sky130_fd_sc_hd__inv_2 _11018_ (.A(\rbzero.map_rom.f1 ),
    .Y(_03746_));
 sky130_fd_sc_hd__o2111a_1 _11019_ (.A1(_03742_),
    .A2(_03743_),
    .B1(_03744_),
    .C1(_03745_),
    .D1(_03746_),
    .X(_03747_));
 sky130_fd_sc_hd__or3_1 _11020_ (.A(\rbzero.map_rom.b6 ),
    .B(\rbzero.map_rom.a6 ),
    .C(\rbzero.map_rom.i_row[4] ),
    .X(_03748_));
 sky130_fd_sc_hd__a211oi_1 _11021_ (.A1(_03738_),
    .A2(_03748_),
    .B1(\rbzero.map_rom.d6 ),
    .C1(\rbzero.map_rom.c6 ),
    .Y(_03749_));
 sky130_fd_sc_hd__a31o_1 _11022_ (.A1(_03740_),
    .A2(_03741_),
    .A3(_03747_),
    .B1(_03749_),
    .X(_03750_));
 sky130_fd_sc_hd__and3_1 _11023_ (.A(_03736_),
    .B(\rbzero.map_rom.f1 ),
    .C(\rbzero.map_rom.i_col[4] ),
    .X(_03751_));
 sky130_fd_sc_hd__or3_1 _11024_ (.A(\rbzero.map_rom.f4 ),
    .B(\rbzero.map_rom.f3 ),
    .C(\rbzero.map_rom.i_col[4] ),
    .X(_03752_));
 sky130_fd_sc_hd__or3_1 _11025_ (.A(_03736_),
    .B(\rbzero.map_rom.f1 ),
    .C(_03752_),
    .X(_03753_));
 sky130_fd_sc_hd__o31ai_1 _11026_ (.A1(\rbzero.map_rom.f4 ),
    .A2(\rbzero.map_rom.d6 ),
    .A3(_03740_),
    .B1(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__a31o_1 _11027_ (.A1(\rbzero.map_rom.f4 ),
    .A2(\rbzero.map_rom.f3 ),
    .A3(_03751_),
    .B1(_03754_),
    .X(_03755_));
 sky130_fd_sc_hd__a311o_1 _11028_ (.A1(\rbzero.map_rom.d6 ),
    .A2(\rbzero.map_rom.c6 ),
    .A3(_03739_),
    .B1(_03750_),
    .C1(_03755_),
    .X(_03756_));
 sky130_fd_sc_hd__xor2_1 _11029_ (.A(_03736_),
    .B(\rbzero.map_rom.a6 ),
    .X(_03757_));
 sky130_fd_sc_hd__nand2_1 _11030_ (.A(\rbzero.map_rom.f1 ),
    .B(\rbzero.map_rom.c6 ),
    .Y(_03758_));
 sky130_fd_sc_hd__o2bb2a_1 _11031_ (.A1_N(\rbzero.map_rom.f4 ),
    .A2_N(_03733_),
    .B1(\rbzero.map_rom.d6 ),
    .B2(\rbzero.map_rom.f3 ),
    .X(_03759_));
 sky130_fd_sc_hd__o211a_1 _11032_ (.A1(\rbzero.map_rom.f4 ),
    .A2(_03733_),
    .B1(_03758_),
    .C1(_03759_),
    .X(_03760_));
 sky130_fd_sc_hd__o221a_1 _11033_ (.A1(_03735_),
    .A2(_03743_),
    .B1(\rbzero.map_rom.c6 ),
    .B2(\rbzero.map_rom.f1 ),
    .C1(_03760_),
    .X(_03761_));
 sky130_fd_sc_hd__or4_1 _11034_ (.A(\rbzero.map_rom.d6 ),
    .B(_03744_),
    .C(\rbzero.map_rom.i_row[4] ),
    .D(_03758_),
    .X(_03762_));
 sky130_fd_sc_hd__or4_1 _11035_ (.A(_03736_),
    .B(_03733_),
    .C(_03752_),
    .D(_03762_),
    .X(_03763_));
 sky130_fd_sc_hd__a21bo_1 _11036_ (.A1(_03757_),
    .A2(_03761_),
    .B1_N(_03763_),
    .X(_03764_));
 sky130_fd_sc_hd__a22o_1 _11037_ (.A1(\rbzero.otherx[0] ),
    .A2(_03742_),
    .B1(_03746_),
    .B2(\rbzero.otherx[3] ),
    .X(_03765_));
 sky130_fd_sc_hd__inv_2 _11038_ (.A(\rbzero.othery[4] ),
    .Y(_03766_));
 sky130_fd_sc_hd__o2bb2a_1 _11039_ (.A1_N(\rbzero.otherx[1] ),
    .A2_N(_03735_),
    .B1(_03746_),
    .B2(\rbzero.otherx[3] ),
    .X(_03767_));
 sky130_fd_sc_hd__o221a_1 _11040_ (.A1(\rbzero.otherx[1] ),
    .A2(_03735_),
    .B1(\rbzero.map_rom.i_row[4] ),
    .B2(_03766_),
    .C1(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__xor2_1 _11041_ (.A(\rbzero.othery[1] ),
    .B(\rbzero.map_rom.c6 ),
    .X(_03769_));
 sky130_fd_sc_hd__xor2_1 _11042_ (.A(\rbzero.otherx[2] ),
    .B(_03736_),
    .X(_03770_));
 sky130_fd_sc_hd__a221o_1 _11043_ (.A1(\rbzero.othery[3] ),
    .A2(_03744_),
    .B1(\rbzero.map_rom.i_row[4] ),
    .B2(_03766_),
    .C1(_03770_),
    .X(_03771_));
 sky130_fd_sc_hd__xnor2_1 _11044_ (.A(\rbzero.othery[2] ),
    .B(_03733_),
    .Y(_03772_));
 sky130_fd_sc_hd__xnor2_1 _11045_ (.A(\rbzero.othery[0] ),
    .B(\rbzero.map_rom.d6 ),
    .Y(_03773_));
 sky130_fd_sc_hd__o221a_1 _11046_ (.A1(\rbzero.otherx[0] ),
    .A2(_03742_),
    .B1(_03744_),
    .B2(\rbzero.othery[3] ),
    .C1(_03773_),
    .X(_03774_));
 sky130_fd_sc_hd__and4bb_1 _11047_ (.A_N(_03769_),
    .B_N(_03771_),
    .C(_03772_),
    .D(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__xnor2_1 _11048_ (.A(\rbzero.otherx[4] ),
    .B(\rbzero.map_rom.i_col[4] ),
    .Y(_03776_));
 sky130_fd_sc_hd__and4b_1 _11049_ (.A_N(_03765_),
    .B(_03768_),
    .C(_03775_),
    .D(_03776_),
    .X(_03777_));
 sky130_fd_sc_hd__nor3_2 _11050_ (.A(_03756_),
    .B(_03764_),
    .C(_03777_),
    .Y(_03778_));
 sky130_fd_sc_hd__or2_1 _11051_ (.A(_03731_),
    .B(_03778_),
    .X(_03779_));
 sky130_fd_sc_hd__nor2_1 _11052_ (.A(_03730_),
    .B(_03779_),
    .Y(_00016_));
 sky130_fd_sc_hd__buf_2 _11053_ (.A(\gpout0.hpos[5] ),
    .X(_03780_));
 sky130_fd_sc_hd__buf_2 _11054_ (.A(_03780_),
    .X(_03781_));
 sky130_fd_sc_hd__and2_1 _11055_ (.A(\gpout0.hpos[3] ),
    .B(\gpout0.hpos[4] ),
    .X(_03782_));
 sky130_fd_sc_hd__clkbuf_4 _11056_ (.A(\gpout0.hpos[6] ),
    .X(_03783_));
 sky130_fd_sc_hd__clkbuf_4 _11057_ (.A(_03783_),
    .X(_03784_));
 sky130_fd_sc_hd__o21ai_1 _11058_ (.A1(_03781_),
    .A2(_03782_),
    .B1(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__or3_1 _11059_ (.A(_03291_),
    .B(_03294_),
    .C(_03296_),
    .X(_03786_));
 sky130_fd_sc_hd__a211o_1 _11060_ (.A1(_03781_),
    .A2(_03782_),
    .B1(_03785_),
    .C1(_03786_),
    .X(_03787_));
 sky130_fd_sc_hd__buf_4 _11061_ (.A(_03787_),
    .X(o_tex_oeb0));
 sky130_fd_sc_hd__inv_2 _11062_ (.A(_03290_),
    .Y(_03788_));
 sky130_fd_sc_hd__a21bo_2 _11063_ (.A1(_03788_),
    .A2(_03785_),
    .B1_N(_03297_),
    .X(o_tex_csb));
 sky130_fd_sc_hd__clkbuf_4 _11064_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_03789_));
 sky130_fd_sc_hd__clkbuf_4 _11065_ (.A(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__inv_2 _11066_ (.A(\rbzero.wall_tracer.state[8] ),
    .Y(_03791_));
 sky130_fd_sc_hd__inv_2 _11067_ (.A(\rbzero.wall_tracer.state[11] ),
    .Y(_03792_));
 sky130_fd_sc_hd__a311o_1 _11068_ (.A1(_03790_),
    .A2(_03791_),
    .A3(_03792_),
    .B1(_03730_),
    .C1(\rbzero.wall_tracer.state[0] ),
    .X(_00011_));
 sky130_fd_sc_hd__clkinv_2 _11069_ (.A(\rbzero.wall_tracer.state[13] ),
    .Y(_03793_));
 sky130_fd_sc_hd__clkbuf_4 _11070_ (.A(_03793_),
    .X(_03794_));
 sky130_fd_sc_hd__buf_4 _11071_ (.A(_03794_),
    .X(_03795_));
 sky130_fd_sc_hd__buf_4 _11072_ (.A(_03795_),
    .X(_03796_));
 sky130_fd_sc_hd__buf_6 _11073_ (.A(\rbzero.wall_tracer.state[1] ),
    .X(_03797_));
 sky130_fd_sc_hd__buf_6 _11074_ (.A(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__nand2_2 _11075_ (.A(_03798_),
    .B(_03778_),
    .Y(_03799_));
 sky130_fd_sc_hd__clkbuf_4 _11076_ (.A(_03799_),
    .X(_03800_));
 sky130_fd_sc_hd__a21oi_1 _11077_ (.A1(_03796_),
    .A2(_03800_),
    .B1(_03730_),
    .Y(_00015_));
 sky130_fd_sc_hd__nor2_1 _11078_ (.A(\rbzero.vga_sync.vsync ),
    .B(_03442_),
    .Y(_03801_));
 sky130_fd_sc_hd__o21ai_2 _11079_ (.A1(_03290_),
    .A2(\gpout0.hpos[8] ),
    .B1(\gpout0.hpos[9] ),
    .Y(_03802_));
 sky130_fd_sc_hd__or2_1 _11080_ (.A(_03783_),
    .B(_03780_),
    .X(_03803_));
 sky130_fd_sc_hd__and3_1 _11081_ (.A(\gpout0.hpos[2] ),
    .B(\gpout0.hpos[1] ),
    .C(\gpout0.hpos[0] ),
    .X(_03804_));
 sky130_fd_sc_hd__and2_1 _11082_ (.A(_03782_),
    .B(_03804_),
    .X(_03805_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11083_ (.A(_03805_),
    .X(_03806_));
 sky130_fd_sc_hd__or3b_2 _11084_ (.A(_03803_),
    .B(_03290_),
    .C_N(_03806_),
    .X(_03807_));
 sky130_fd_sc_hd__nor2_4 _11085_ (.A(_03802_),
    .B(_03807_),
    .Y(_03808_));
 sky130_fd_sc_hd__nand2_4 _11086_ (.A(\rbzero.wall_tracer.state[14] ),
    .B(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__and2_1 _11087_ (.A(_03801_),
    .B(_03809_),
    .X(_03810_));
 sky130_fd_sc_hd__clkinv_2 _11088_ (.A(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__clkbuf_4 _11089_ (.A(_03811_),
    .X(_03812_));
 sky130_fd_sc_hd__buf_4 _11090_ (.A(_03812_),
    .X(_00013_));
 sky130_fd_sc_hd__or2_2 _11091_ (.A(_03802_),
    .B(_03807_),
    .X(_03813_));
 sky130_fd_sc_hd__a21oi_1 _11092_ (.A1(\rbzero.wall_tracer.state[14] ),
    .A2(_03813_),
    .B1(\rbzero.wall_tracer.state[10] ),
    .Y(_03814_));
 sky130_fd_sc_hd__nor2_1 _11093_ (.A(_03730_),
    .B(_03814_),
    .Y(_00014_));
 sky130_fd_sc_hd__nor2_1 _11094_ (.A(_03792_),
    .B(_03729_),
    .Y(_00000_));
 sky130_fd_sc_hd__buf_2 _11095_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_03815_));
 sky130_fd_sc_hd__clkbuf_4 _11096_ (.A(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__inv_2 _11097_ (.A(\rbzero.wall_tracer.state[0] ),
    .Y(_03817_));
 sky130_fd_sc_hd__clkbuf_4 _11098_ (.A(_03801_),
    .X(_03818_));
 sky130_fd_sc_hd__buf_4 _11099_ (.A(_03818_),
    .X(_03819_));
 sky130_fd_sc_hd__a41o_1 _11100_ (.A1(_03816_),
    .A2(_03817_),
    .A3(_03791_),
    .A4(_03819_),
    .B1(_00000_),
    .X(_00012_));
 sky130_fd_sc_hd__or4b_1 _11101_ (.A(\gpout0.vpos[9] ),
    .B(\gpout0.vpos[8] ),
    .C(\gpout0.vpos[7] ),
    .D_N(net2),
    .X(_03820_));
 sky130_fd_sc_hd__or3_2 _11102_ (.A(\gpout0.vpos[5] ),
    .B(\gpout0.vpos[4] ),
    .C(\gpout0.vpos[3] ),
    .X(_03821_));
 sky130_fd_sc_hd__o41a_1 _11103_ (.A1(\gpout0.vpos[2] ),
    .A2(\gpout0.vpos[1] ),
    .A3(\gpout0.vpos[0] ),
    .A4(_03821_),
    .B1(\gpout0.vpos[6] ),
    .X(_03822_));
 sky130_fd_sc_hd__a31o_1 _11104_ (.A1(\gpout0.hpos[5] ),
    .A2(_03782_),
    .A3(_03804_),
    .B1(\gpout0.hpos[6] ),
    .X(_03823_));
 sky130_fd_sc_hd__a31o_1 _11105_ (.A1(\gpout0.hpos[7] ),
    .A2(\gpout0.hpos[8] ),
    .A3(_03823_),
    .B1(\gpout0.hpos[9] ),
    .X(_03824_));
 sky130_fd_sc_hd__or3b_2 _11106_ (.A(_03820_),
    .B(_03822_),
    .C_N(_03824_),
    .X(_03825_));
 sky130_fd_sc_hd__clkinv_2 _11107_ (.A(_03825_),
    .Y(_03826_));
 sky130_fd_sc_hd__nand2_1 _11108_ (.A(\rbzero.traced_texVinit[6] ),
    .B(\rbzero.spi_registers.vshift[3] ),
    .Y(_03827_));
 sky130_fd_sc_hd__or2_1 _11109_ (.A(\rbzero.traced_texVinit[6] ),
    .B(\rbzero.spi_registers.vshift[3] ),
    .X(_03828_));
 sky130_fd_sc_hd__nand3_1 _11110_ (.A(\rbzero.texV[6] ),
    .B(_03827_),
    .C(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__and2_1 _11111_ (.A(\rbzero.traced_texVinit[7] ),
    .B(\rbzero.spi_registers.vshift[4] ),
    .X(_03830_));
 sky130_fd_sc_hd__nor2_1 _11112_ (.A(\rbzero.traced_texVinit[7] ),
    .B(\rbzero.spi_registers.vshift[4] ),
    .Y(_03831_));
 sky130_fd_sc_hd__nor2_1 _11113_ (.A(_03830_),
    .B(_03831_),
    .Y(_03832_));
 sky130_fd_sc_hd__xnor2_1 _11114_ (.A(\rbzero.texV[7] ),
    .B(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__a21oi_1 _11115_ (.A1(_03827_),
    .A2(_03829_),
    .B1(_03833_),
    .Y(_03834_));
 sky130_fd_sc_hd__a21o_1 _11116_ (.A1(_03827_),
    .A2(_03828_),
    .B1(\rbzero.texV[6] ),
    .X(_03835_));
 sky130_fd_sc_hd__nand2_1 _11117_ (.A(_03829_),
    .B(_03835_),
    .Y(_03836_));
 sky130_fd_sc_hd__or2_1 _11118_ (.A(\rbzero.traced_texVinit[5] ),
    .B(\rbzero.spi_registers.vshift[2] ),
    .X(_03837_));
 sky130_fd_sc_hd__nand2_1 _11119_ (.A(\rbzero.traced_texVinit[5] ),
    .B(\rbzero.spi_registers.vshift[2] ),
    .Y(_03838_));
 sky130_fd_sc_hd__a21boi_1 _11120_ (.A1(\rbzero.texV[5] ),
    .A2(_03837_),
    .B1_N(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__nor2_1 _11121_ (.A(_03836_),
    .B(_03839_),
    .Y(_03840_));
 sky130_fd_sc_hd__nand2_1 _11122_ (.A(_03838_),
    .B(_03837_),
    .Y(_03841_));
 sky130_fd_sc_hd__xor2_1 _11123_ (.A(\rbzero.texV[5] ),
    .B(_03841_),
    .X(_03842_));
 sky130_fd_sc_hd__or2_1 _11124_ (.A(\rbzero.traced_texVinit[4] ),
    .B(\rbzero.spi_registers.vshift[1] ),
    .X(_03843_));
 sky130_fd_sc_hd__nand2_1 _11125_ (.A(\rbzero.traced_texVinit[4] ),
    .B(\rbzero.spi_registers.vshift[1] ),
    .Y(_03844_));
 sky130_fd_sc_hd__a21boi_1 _11126_ (.A1(\rbzero.texV[4] ),
    .A2(_03843_),
    .B1_N(_03844_),
    .Y(_03845_));
 sky130_fd_sc_hd__nor2_1 _11127_ (.A(_03842_),
    .B(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__nand2_1 _11128_ (.A(_03844_),
    .B(_03843_),
    .Y(_03847_));
 sky130_fd_sc_hd__xor2_1 _11129_ (.A(\rbzero.texV[4] ),
    .B(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__or2_1 _11130_ (.A(\rbzero.traced_texVinit[3] ),
    .B(\rbzero.spi_registers.vshift[0] ),
    .X(_03849_));
 sky130_fd_sc_hd__nand2_1 _11131_ (.A(\rbzero.traced_texVinit[3] ),
    .B(\rbzero.spi_registers.vshift[0] ),
    .Y(_03850_));
 sky130_fd_sc_hd__a21boi_1 _11132_ (.A1(\rbzero.texV[3] ),
    .A2(_03849_),
    .B1_N(_03850_),
    .Y(_03851_));
 sky130_fd_sc_hd__nor2_1 _11133_ (.A(_03848_),
    .B(_03851_),
    .Y(_03852_));
 sky130_fd_sc_hd__xnor2_1 _11134_ (.A(_03848_),
    .B(_03851_),
    .Y(_03853_));
 sky130_fd_sc_hd__nand2_1 _11135_ (.A(_03850_),
    .B(_03849_),
    .Y(_03854_));
 sky130_fd_sc_hd__xor2_1 _11136_ (.A(\rbzero.texV[3] ),
    .B(_03854_),
    .X(_03855_));
 sky130_fd_sc_hd__o211a_1 _11137_ (.A1(\rbzero.traced_texVinit[1] ),
    .A2(\rbzero.texV[1] ),
    .B1(\rbzero.texV[0] ),
    .C1(\rbzero.traced_texVinit[0] ),
    .X(_03856_));
 sky130_fd_sc_hd__a221o_1 _11138_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(\rbzero.texV[2] ),
    .B1(\rbzero.texV[1] ),
    .B2(\rbzero.traced_texVinit[1] ),
    .C1(_03856_),
    .X(_03857_));
 sky130_fd_sc_hd__o21ai_2 _11139_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(\rbzero.texV[2] ),
    .B1(_03857_),
    .Y(_03858_));
 sky130_fd_sc_hd__or2_2 _11140_ (.A(_03855_),
    .B(_03858_),
    .X(_03859_));
 sky130_fd_sc_hd__nor2_2 _11141_ (.A(_03853_),
    .B(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hd__and2_1 _11142_ (.A(_03842_),
    .B(_03845_),
    .X(_03861_));
 sky130_fd_sc_hd__or2_1 _11143_ (.A(_03846_),
    .B(_03861_),
    .X(_03862_));
 sky130_fd_sc_hd__inv_2 _11144_ (.A(_03862_),
    .Y(_03863_));
 sky130_fd_sc_hd__o21a_1 _11145_ (.A1(_03852_),
    .A2(_03860_),
    .B1(_03863_),
    .X(_03864_));
 sky130_fd_sc_hd__and2_1 _11146_ (.A(_03836_),
    .B(_03839_),
    .X(_03865_));
 sky130_fd_sc_hd__or2_1 _11147_ (.A(_03840_),
    .B(_03865_),
    .X(_03866_));
 sky130_fd_sc_hd__inv_2 _11148_ (.A(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__o21a_1 _11149_ (.A1(_03846_),
    .A2(_03864_),
    .B1(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__and3_1 _11150_ (.A(_03833_),
    .B(_03827_),
    .C(_03829_),
    .X(_03869_));
 sky130_fd_sc_hd__or2_1 _11151_ (.A(_03834_),
    .B(_03869_),
    .X(_03870_));
 sky130_fd_sc_hd__inv_2 _11152_ (.A(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__o21a_1 _11153_ (.A1(_03840_),
    .A2(_03868_),
    .B1(_03871_),
    .X(_03872_));
 sky130_fd_sc_hd__and2_1 _11154_ (.A(\rbzero.traced_texVinit[8] ),
    .B(\rbzero.spi_registers.vshift[5] ),
    .X(_03873_));
 sky130_fd_sc_hd__nor2_1 _11155_ (.A(\rbzero.traced_texVinit[8] ),
    .B(\rbzero.spi_registers.vshift[5] ),
    .Y(_03874_));
 sky130_fd_sc_hd__nor2_1 _11156_ (.A(_03873_),
    .B(_03874_),
    .Y(_03875_));
 sky130_fd_sc_hd__xnor2_1 _11157_ (.A(\rbzero.texV[8] ),
    .B(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hd__a21oi_1 _11158_ (.A1(\rbzero.texV[7] ),
    .A2(_03832_),
    .B1(_03830_),
    .Y(_03877_));
 sky130_fd_sc_hd__xnor2_1 _11159_ (.A(_03876_),
    .B(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__o21ba_2 _11160_ (.A1(_03834_),
    .A2(_03872_),
    .B1_N(_03878_),
    .X(_03879_));
 sky130_fd_sc_hd__nand2_1 _11161_ (.A(\rbzero.traced_texVinit[10] ),
    .B(\rbzero.texV[10] ),
    .Y(_03880_));
 sky130_fd_sc_hd__or2_1 _11162_ (.A(\rbzero.traced_texVinit[10] ),
    .B(\rbzero.texV[10] ),
    .X(_03881_));
 sky130_fd_sc_hd__xnor2_1 _11163_ (.A(\rbzero.traced_texVinit[9] ),
    .B(\rbzero.texV[9] ),
    .Y(_03882_));
 sky130_fd_sc_hd__a21oi_1 _11164_ (.A1(\rbzero.texV[8] ),
    .A2(_03875_),
    .B1(_03873_),
    .Y(_03883_));
 sky130_fd_sc_hd__o22ai_1 _11165_ (.A1(_03876_),
    .A2(_03877_),
    .B1(_03882_),
    .B2(_03883_),
    .Y(_03884_));
 sky130_fd_sc_hd__a22o_1 _11166_ (.A1(\rbzero.traced_texVinit[9] ),
    .A2(\rbzero.texV[9] ),
    .B1(_03880_),
    .B2(_03881_),
    .X(_03885_));
 sky130_fd_sc_hd__nand2_1 _11167_ (.A(_03882_),
    .B(_03883_),
    .Y(_03886_));
 sky130_fd_sc_hd__o211a_1 _11168_ (.A1(_03879_),
    .A2(_03884_),
    .B1(_03885_),
    .C1(_03886_),
    .X(_03887_));
 sky130_fd_sc_hd__a41o_1 _11169_ (.A1(\rbzero.traced_texVinit[9] ),
    .A2(\rbzero.texV[9] ),
    .A3(_03880_),
    .A4(_03881_),
    .B1(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__xnor2_1 _11170_ (.A(\rbzero.traced_texVinit[11] ),
    .B(\rbzero.texV[11] ),
    .Y(_03889_));
 sky130_fd_sc_hd__xnor2_1 _11171_ (.A(_03880_),
    .B(_03889_),
    .Y(_03890_));
 sky130_fd_sc_hd__nand2_1 _11172_ (.A(_03888_),
    .B(_03890_),
    .Y(_03891_));
 sky130_fd_sc_hd__or2_1 _11173_ (.A(_03888_),
    .B(_03890_),
    .X(_03892_));
 sky130_fd_sc_hd__a21oi_1 _11174_ (.A1(_03891_),
    .A2(_03892_),
    .B1(\rbzero.row_render.vinf ),
    .Y(_03893_));
 sky130_fd_sc_hd__buf_4 _11175_ (.A(_03893_),
    .X(_03894_));
 sky130_fd_sc_hd__nor3b_2 _11176_ (.A(_03834_),
    .B(_03872_),
    .C_N(_03878_),
    .Y(_03895_));
 sky130_fd_sc_hd__or3_4 _11177_ (.A(_03879_),
    .B(_03894_),
    .C(_03895_),
    .X(_03896_));
 sky130_fd_sc_hd__nor3_1 _11178_ (.A(_03867_),
    .B(_03846_),
    .C(_03864_),
    .Y(_03897_));
 sky130_fd_sc_hd__nor3_4 _11179_ (.A(_03868_),
    .B(_03894_),
    .C(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__buf_4 _11180_ (.A(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__buf_4 _11181_ (.A(_03899_),
    .X(_03900_));
 sky130_fd_sc_hd__a21oi_2 _11182_ (.A1(_03855_),
    .A2(_03858_),
    .B1(_03893_),
    .Y(_03901_));
 sky130_fd_sc_hd__nand2_1 _11183_ (.A(_03859_),
    .B(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__buf_2 _11184_ (.A(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__buf_4 _11185_ (.A(_03903_),
    .X(_03904_));
 sky130_fd_sc_hd__mux2_1 _11186_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_03904_),
    .X(_03905_));
 sky130_fd_sc_hd__mux2_1 _11187_ (.A0(\rbzero.tex_r0[51] ),
    .A1(\rbzero.tex_r0[50] ),
    .S(_03904_),
    .X(_03906_));
 sky130_fd_sc_hd__nand2_1 _11188_ (.A(_03853_),
    .B(_03859_),
    .Y(_03907_));
 sky130_fd_sc_hd__nor3b_4 _11189_ (.A(_03860_),
    .B(_03894_),
    .C_N(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__buf_4 _11190_ (.A(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__buf_4 _11191_ (.A(_03909_),
    .X(_03910_));
 sky130_fd_sc_hd__mux2_1 _11192_ (.A0(_03905_),
    .A1(_03906_),
    .S(_03910_),
    .X(_03911_));
 sky130_fd_sc_hd__mux2_1 _11193_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(_03904_),
    .X(_03912_));
 sky130_fd_sc_hd__mux2_1 _11194_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(_03904_),
    .X(_03913_));
 sky130_fd_sc_hd__or3b_2 _11195_ (.A(_03860_),
    .B(_03894_),
    .C_N(_03907_),
    .X(_03914_));
 sky130_fd_sc_hd__buf_4 _11196_ (.A(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__buf_6 _11197_ (.A(_03915_),
    .X(_03916_));
 sky130_fd_sc_hd__mux2_1 _11198_ (.A0(_03912_),
    .A1(_03913_),
    .S(_03916_),
    .X(_03917_));
 sky130_fd_sc_hd__nor3_1 _11199_ (.A(_03863_),
    .B(_03852_),
    .C(_03860_),
    .Y(_03918_));
 sky130_fd_sc_hd__nor3_2 _11200_ (.A(_03864_),
    .B(_03894_),
    .C(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__clkbuf_4 _11201_ (.A(_03919_),
    .X(_03920_));
 sky130_fd_sc_hd__buf_4 _11202_ (.A(_03920_),
    .X(_03921_));
 sky130_fd_sc_hd__mux2_1 _11203_ (.A0(_03911_),
    .A1(_03917_),
    .S(_03921_),
    .X(_03922_));
 sky130_fd_sc_hd__buf_4 _11204_ (.A(_03920_),
    .X(_03923_));
 sky130_fd_sc_hd__buf_4 _11205_ (.A(_03923_),
    .X(_03924_));
 sky130_fd_sc_hd__buf_4 _11206_ (.A(_03903_),
    .X(_03925_));
 sky130_fd_sc_hd__mux2_1 _11207_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_03925_),
    .X(_03926_));
 sky130_fd_sc_hd__mux2_1 _11208_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_03925_),
    .X(_03927_));
 sky130_fd_sc_hd__clkbuf_4 _11209_ (.A(_03914_),
    .X(_03928_));
 sky130_fd_sc_hd__buf_4 _11210_ (.A(_03928_),
    .X(_03929_));
 sky130_fd_sc_hd__buf_4 _11211_ (.A(_03929_),
    .X(_03930_));
 sky130_fd_sc_hd__mux2_1 _11212_ (.A0(_03926_),
    .A1(_03927_),
    .S(_03930_),
    .X(_03931_));
 sky130_fd_sc_hd__clkbuf_4 _11213_ (.A(_03909_),
    .X(_03932_));
 sky130_fd_sc_hd__mux2_1 _11214_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(_03925_),
    .X(_03933_));
 sky130_fd_sc_hd__clkbuf_4 _11215_ (.A(_03902_),
    .X(_03934_));
 sky130_fd_sc_hd__buf_4 _11216_ (.A(_03934_),
    .X(_03935_));
 sky130_fd_sc_hd__buf_4 _11217_ (.A(_03935_),
    .X(_03936_));
 sky130_fd_sc_hd__and2_1 _11218_ (.A(\rbzero.tex_r0[58] ),
    .B(_03936_),
    .X(_03937_));
 sky130_fd_sc_hd__clkbuf_4 _11219_ (.A(_03859_),
    .X(_03938_));
 sky130_fd_sc_hd__clkbuf_4 _11220_ (.A(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__clkbuf_4 _11221_ (.A(_03901_),
    .X(_03940_));
 sky130_fd_sc_hd__clkbuf_4 _11222_ (.A(_03940_),
    .X(_03941_));
 sky130_fd_sc_hd__buf_4 _11223_ (.A(_03915_),
    .X(_03942_));
 sky130_fd_sc_hd__a31o_1 _11224_ (.A1(\rbzero.tex_r0[59] ),
    .A2(_03939_),
    .A3(_03941_),
    .B1(_03942_),
    .X(_03943_));
 sky130_fd_sc_hd__or3_4 _11225_ (.A(_03864_),
    .B(_03894_),
    .C(_03918_),
    .X(_03944_));
 sky130_fd_sc_hd__buf_4 _11226_ (.A(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__clkbuf_4 _11227_ (.A(_03945_),
    .X(_03946_));
 sky130_fd_sc_hd__o221a_1 _11228_ (.A1(_03932_),
    .A2(_03933_),
    .B1(_03937_),
    .B2(_03943_),
    .C1(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__or3_1 _11229_ (.A(_03868_),
    .B(_03894_),
    .C(_03897_),
    .X(_03948_));
 sky130_fd_sc_hd__clkbuf_4 _11230_ (.A(_03948_),
    .X(_03949_));
 sky130_fd_sc_hd__clkbuf_4 _11231_ (.A(_03949_),
    .X(_03950_));
 sky130_fd_sc_hd__a211o_1 _11232_ (.A1(_03924_),
    .A2(_03931_),
    .B1(_03947_),
    .C1(_03950_),
    .X(_03951_));
 sky130_fd_sc_hd__nor3_1 _11233_ (.A(_03871_),
    .B(_03840_),
    .C(_03868_),
    .Y(_03952_));
 sky130_fd_sc_hd__nor3_2 _11234_ (.A(_03872_),
    .B(_03894_),
    .C(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__buf_4 _11235_ (.A(_03953_),
    .X(_03954_));
 sky130_fd_sc_hd__o211a_1 _11236_ (.A1(_03900_),
    .A2(_03922_),
    .B1(_03951_),
    .C1(_03954_),
    .X(_03955_));
 sky130_fd_sc_hd__buf_4 _11237_ (.A(_03949_),
    .X(_03956_));
 sky130_fd_sc_hd__buf_4 _11238_ (.A(_03909_),
    .X(_03957_));
 sky130_fd_sc_hd__clkbuf_4 _11239_ (.A(_03957_),
    .X(_03958_));
 sky130_fd_sc_hd__clkbuf_4 _11240_ (.A(_03925_),
    .X(_03959_));
 sky130_fd_sc_hd__mux2_1 _11241_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_03959_),
    .X(_03960_));
 sky130_fd_sc_hd__buf_4 _11242_ (.A(_03903_),
    .X(_03961_));
 sky130_fd_sc_hd__clkbuf_4 _11243_ (.A(_03961_),
    .X(_03962_));
 sky130_fd_sc_hd__and2_1 _11244_ (.A(\rbzero.tex_r0[46] ),
    .B(_03962_),
    .X(_03963_));
 sky130_fd_sc_hd__buf_2 _11245_ (.A(_03939_),
    .X(_03964_));
 sky130_fd_sc_hd__clkbuf_4 _11246_ (.A(_03941_),
    .X(_03965_));
 sky130_fd_sc_hd__a31o_1 _11247_ (.A1(\rbzero.tex_r0[47] ),
    .A2(_03964_),
    .A3(_03965_),
    .B1(_03930_),
    .X(_03966_));
 sky130_fd_sc_hd__o221a_1 _11248_ (.A1(_03958_),
    .A2(_03960_),
    .B1(_03963_),
    .B2(_03966_),
    .C1(_03924_),
    .X(_03967_));
 sky130_fd_sc_hd__buf_4 _11249_ (.A(_03916_),
    .X(_03968_));
 sky130_fd_sc_hd__mux2_1 _11250_ (.A0(\rbzero.tex_r0[43] ),
    .A1(\rbzero.tex_r0[42] ),
    .S(_03959_),
    .X(_03969_));
 sky130_fd_sc_hd__and2_1 _11251_ (.A(\rbzero.tex_r0[40] ),
    .B(_03962_),
    .X(_03970_));
 sky130_fd_sc_hd__a31o_1 _11252_ (.A1(\rbzero.tex_r0[41] ),
    .A2(_03964_),
    .A3(_03965_),
    .B1(_03932_),
    .X(_03971_));
 sky130_fd_sc_hd__buf_4 _11253_ (.A(_03945_),
    .X(_03972_));
 sky130_fd_sc_hd__o221a_1 _11254_ (.A1(_03968_),
    .A2(_03969_),
    .B1(_03970_),
    .B2(_03971_),
    .C1(_03972_),
    .X(_03973_));
 sky130_fd_sc_hd__buf_4 _11255_ (.A(_03903_),
    .X(_03974_));
 sky130_fd_sc_hd__mux2_1 _11256_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_03974_),
    .X(_03975_));
 sky130_fd_sc_hd__mux2_1 _11257_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_03974_),
    .X(_03976_));
 sky130_fd_sc_hd__mux2_1 _11258_ (.A0(_03975_),
    .A1(_03976_),
    .S(_03930_),
    .X(_03977_));
 sky130_fd_sc_hd__mux2_1 _11259_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_03974_),
    .X(_03978_));
 sky130_fd_sc_hd__and3_1 _11260_ (.A(\rbzero.tex_r0[35] ),
    .B(_03939_),
    .C(_03941_),
    .X(_03979_));
 sky130_fd_sc_hd__buf_4 _11261_ (.A(_03935_),
    .X(_03980_));
 sky130_fd_sc_hd__a21o_1 _11262_ (.A1(\rbzero.tex_r0[34] ),
    .A2(_03980_),
    .B1(_03942_),
    .X(_03981_));
 sky130_fd_sc_hd__o221a_1 _11263_ (.A1(_03932_),
    .A2(_03978_),
    .B1(_03979_),
    .B2(_03981_),
    .C1(_03946_),
    .X(_03982_));
 sky130_fd_sc_hd__a211o_1 _11264_ (.A1(_03924_),
    .A2(_03977_),
    .B1(_03982_),
    .C1(_03899_),
    .X(_03983_));
 sky130_fd_sc_hd__or3_2 _11265_ (.A(_03872_),
    .B(_03894_),
    .C(_03952_),
    .X(_03984_));
 sky130_fd_sc_hd__buf_6 _11266_ (.A(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__o311a_1 _11267_ (.A1(_03956_),
    .A2(_03967_),
    .A3(_03973_),
    .B1(_03983_),
    .C1(_03985_),
    .X(_03986_));
 sky130_fd_sc_hd__mux2_1 _11268_ (.A0(\rbzero.tex_r0[19] ),
    .A1(\rbzero.tex_r0[18] ),
    .S(_03974_),
    .X(_03987_));
 sky130_fd_sc_hd__mux2_1 _11269_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_03974_),
    .X(_03988_));
 sky130_fd_sc_hd__mux2_1 _11270_ (.A0(_03987_),
    .A1(_03988_),
    .S(_03930_),
    .X(_03989_));
 sky130_fd_sc_hd__mux2_1 _11271_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(_03974_),
    .X(_03990_));
 sky130_fd_sc_hd__mux2_1 _11272_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(_03974_),
    .X(_03991_));
 sky130_fd_sc_hd__mux2_1 _11273_ (.A0(_03990_),
    .A1(_03991_),
    .S(_03957_),
    .X(_03992_));
 sky130_fd_sc_hd__mux2_1 _11274_ (.A0(_03989_),
    .A1(_03992_),
    .S(_03924_),
    .X(_03993_));
 sky130_fd_sc_hd__clkbuf_4 _11275_ (.A(_03946_),
    .X(_03994_));
 sky130_fd_sc_hd__mux2_1 _11276_ (.A0(\rbzero.tex_r0[27] ),
    .A1(\rbzero.tex_r0[26] ),
    .S(_03936_),
    .X(_03995_));
 sky130_fd_sc_hd__mux2_1 _11277_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_03936_),
    .X(_03996_));
 sky130_fd_sc_hd__clkbuf_4 _11278_ (.A(_03942_),
    .X(_03997_));
 sky130_fd_sc_hd__mux2_1 _11279_ (.A0(_03995_),
    .A1(_03996_),
    .S(_03997_),
    .X(_03998_));
 sky130_fd_sc_hd__mux2_1 _11280_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_03936_),
    .X(_03999_));
 sky130_fd_sc_hd__buf_4 _11281_ (.A(_03903_),
    .X(_04000_));
 sky130_fd_sc_hd__buf_4 _11282_ (.A(_04000_),
    .X(_04001_));
 sky130_fd_sc_hd__and2_1 _11283_ (.A(\rbzero.tex_r0[30] ),
    .B(_04001_),
    .X(_04002_));
 sky130_fd_sc_hd__a31o_1 _11284_ (.A1(\rbzero.tex_r0[31] ),
    .A2(_03939_),
    .A3(_03941_),
    .B1(_03942_),
    .X(_04003_));
 sky130_fd_sc_hd__o221a_1 _11285_ (.A1(_03932_),
    .A2(_03999_),
    .B1(_04002_),
    .B2(_04003_),
    .C1(_03923_),
    .X(_04004_));
 sky130_fd_sc_hd__a211o_1 _11286_ (.A1(_03994_),
    .A2(_03998_),
    .B1(_04004_),
    .C1(_03956_),
    .X(_04005_));
 sky130_fd_sc_hd__o211a_1 _11287_ (.A1(_03900_),
    .A2(_03993_),
    .B1(_04005_),
    .C1(_03954_),
    .X(_04006_));
 sky130_fd_sc_hd__buf_4 _11288_ (.A(_03923_),
    .X(_04007_));
 sky130_fd_sc_hd__mux2_1 _11289_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(_03961_),
    .X(_04008_));
 sky130_fd_sc_hd__mux2_1 _11290_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(_03961_),
    .X(_04009_));
 sky130_fd_sc_hd__mux2_1 _11291_ (.A0(_04008_),
    .A1(_04009_),
    .S(_03930_),
    .X(_04010_));
 sky130_fd_sc_hd__mux2_1 _11292_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_03961_),
    .X(_04011_));
 sky130_fd_sc_hd__and3_1 _11293_ (.A(\rbzero.tex_r0[11] ),
    .B(_03939_),
    .C(_03941_),
    .X(_04012_));
 sky130_fd_sc_hd__buf_4 _11294_ (.A(_03904_),
    .X(_04013_));
 sky130_fd_sc_hd__buf_4 _11295_ (.A(_03915_),
    .X(_04014_));
 sky130_fd_sc_hd__a21o_1 _11296_ (.A1(\rbzero.tex_r0[10] ),
    .A2(_04013_),
    .B1(_04014_),
    .X(_04015_));
 sky130_fd_sc_hd__o221a_1 _11297_ (.A1(_03932_),
    .A2(_04011_),
    .B1(_04012_),
    .B2(_04015_),
    .C1(_03946_),
    .X(_04016_));
 sky130_fd_sc_hd__a211o_1 _11298_ (.A1(_04007_),
    .A2(_04010_),
    .B1(_04016_),
    .C1(_03950_),
    .X(_04017_));
 sky130_fd_sc_hd__mux2_1 _11299_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_03961_),
    .X(_04018_));
 sky130_fd_sc_hd__mux2_1 _11300_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_03961_),
    .X(_04019_));
 sky130_fd_sc_hd__mux2_1 _11301_ (.A0(_04018_),
    .A1(_04019_),
    .S(_03932_),
    .X(_04020_));
 sky130_fd_sc_hd__and3_1 _11302_ (.A(\rbzero.tex_r0[3] ),
    .B(_03939_),
    .C(_03941_),
    .X(_04021_));
 sky130_fd_sc_hd__a21o_1 _11303_ (.A1(\rbzero.tex_r0[2] ),
    .A2(_04001_),
    .B1(_03942_),
    .X(_04022_));
 sky130_fd_sc_hd__mux2_1 _11304_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_03936_),
    .X(_04023_));
 sky130_fd_sc_hd__o221a_1 _11305_ (.A1(_04021_),
    .A2(_04022_),
    .B1(_04023_),
    .B2(_03932_),
    .C1(_03946_),
    .X(_04024_));
 sky130_fd_sc_hd__a211o_1 _11306_ (.A1(_04007_),
    .A2(_04020_),
    .B1(_04024_),
    .C1(_03899_),
    .X(_04025_));
 sky130_fd_sc_hd__nor3_4 _11307_ (.A(_03879_),
    .B(_03894_),
    .C(_03895_),
    .Y(_04026_));
 sky130_fd_sc_hd__a31o_1 _11308_ (.A1(_03985_),
    .A2(_04017_),
    .A3(_04025_),
    .B1(_04026_),
    .X(_04027_));
 sky130_fd_sc_hd__o32a_1 _11309_ (.A1(_03896_),
    .A2(_03955_),
    .A3(_03986_),
    .B1(_04006_),
    .B2(_04027_),
    .X(_04028_));
 sky130_fd_sc_hd__o21a_1 _11310_ (.A1(_03784_),
    .A2(_03290_),
    .B1(_03293_),
    .X(_04029_));
 sky130_fd_sc_hd__nor2_4 _11311_ (.A(\gpout0.hpos[9] ),
    .B(_04029_),
    .Y(_04030_));
 sky130_fd_sc_hd__mux2_1 _11312_ (.A0(\rbzero.color_sky[0] ),
    .A1(\rbzero.color_floor[0] ),
    .S(_04030_),
    .X(_04031_));
 sky130_fd_sc_hd__buf_4 _11313_ (.A(_03902_),
    .X(_04032_));
 sky130_fd_sc_hd__o211a_1 _11314_ (.A1(\rbzero.floor_leak[1] ),
    .A2(_03914_),
    .B1(_04032_),
    .C1(\rbzero.floor_leak[0] ),
    .X(_04033_));
 sky130_fd_sc_hd__a221o_1 _11315_ (.A1(\rbzero.floor_leak[1] ),
    .A2(_03928_),
    .B1(_03944_),
    .B2(\rbzero.floor_leak[2] ),
    .C1(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__o221a_1 _11316_ (.A1(\rbzero.floor_leak[2] ),
    .A2(_03945_),
    .B1(_03949_),
    .B2(\rbzero.floor_leak[3] ),
    .C1(_04034_),
    .X(_04035_));
 sky130_fd_sc_hd__a221o_1 _11317_ (.A1(\rbzero.floor_leak[3] ),
    .A2(_03949_),
    .B1(_03984_),
    .B2(\rbzero.floor_leak[4] ),
    .C1(_04035_),
    .X(_04036_));
 sky130_fd_sc_hd__o22a_1 _11318_ (.A1(\rbzero.floor_leak[5] ),
    .A2(_03896_),
    .B1(_03984_),
    .B2(\rbzero.floor_leak[4] ),
    .X(_04037_));
 sky130_fd_sc_hd__and2_1 _11319_ (.A(_03938_),
    .B(_03940_),
    .X(_04038_));
 sky130_fd_sc_hd__or4_1 _11320_ (.A(_04026_),
    .B(_03908_),
    .C(_03898_),
    .D(_04030_),
    .X(_04039_));
 sky130_fd_sc_hd__or4_1 _11321_ (.A(_04038_),
    .B(_03919_),
    .C(_03953_),
    .D(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__inv_2 _11322_ (.A(\rbzero.row_render.size[2] ),
    .Y(_04041_));
 sky130_fd_sc_hd__nor2_1 _11323_ (.A(\rbzero.row_render.size[1] ),
    .B(\rbzero.row_render.size[0] ),
    .Y(_04042_));
 sky130_fd_sc_hd__nand2_1 _11324_ (.A(_04041_),
    .B(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__or2_1 _11325_ (.A(\rbzero.row_render.size[3] ),
    .B(_04043_),
    .X(_04044_));
 sky130_fd_sc_hd__or3_1 _11326_ (.A(\rbzero.row_render.size[5] ),
    .B(\rbzero.row_render.size[4] ),
    .C(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__and2_1 _11327_ (.A(\rbzero.row_render.size[6] ),
    .B(_04045_),
    .X(_04046_));
 sky130_fd_sc_hd__o21a_1 _11328_ (.A1(\rbzero.row_render.size[7] ),
    .A2(_04046_),
    .B1(\rbzero.row_render.size[8] ),
    .X(_04047_));
 sky130_fd_sc_hd__a21o_1 _11329_ (.A1(\rbzero.row_render.size[7] ),
    .A2(\rbzero.row_render.size[6] ),
    .B1(\rbzero.row_render.size[8] ),
    .X(_04048_));
 sky130_fd_sc_hd__nand3_1 _11330_ (.A(\rbzero.row_render.size[8] ),
    .B(\rbzero.row_render.size[7] ),
    .C(\rbzero.row_render.size[6] ),
    .Y(_04049_));
 sky130_fd_sc_hd__and2_1 _11331_ (.A(_04048_),
    .B(_04049_),
    .X(_04050_));
 sky130_fd_sc_hd__nor2_1 _11332_ (.A(\rbzero.row_render.size[9] ),
    .B(_04048_),
    .Y(_04051_));
 sky130_fd_sc_hd__xnor2_1 _11333_ (.A(\rbzero.row_render.size[7] ),
    .B(\rbzero.row_render.size[6] ),
    .Y(_04052_));
 sky130_fd_sc_hd__inv_2 _11334_ (.A(\rbzero.row_render.size[5] ),
    .Y(_04053_));
 sky130_fd_sc_hd__inv_2 _11335_ (.A(\rbzero.row_render.size[4] ),
    .Y(_04054_));
 sky130_fd_sc_hd__inv_2 _11336_ (.A(\rbzero.row_render.size[3] ),
    .Y(_04055_));
 sky130_fd_sc_hd__inv_2 _11337_ (.A(\rbzero.row_render.size[1] ),
    .Y(_04056_));
 sky130_fd_sc_hd__inv_2 _11338_ (.A(\rbzero.row_render.size[0] ),
    .Y(_04057_));
 sky130_fd_sc_hd__o211a_1 _11339_ (.A1(_04056_),
    .A2(\gpout0.hpos[1] ),
    .B1(\gpout0.hpos[0] ),
    .C1(_04057_),
    .X(_04058_));
 sky130_fd_sc_hd__a221o_1 _11340_ (.A1(_04041_),
    .A2(\gpout0.hpos[2] ),
    .B1(\gpout0.hpos[1] ),
    .B2(_04056_),
    .C1(_04058_),
    .X(_04059_));
 sky130_fd_sc_hd__o221a_1 _11341_ (.A1(_04055_),
    .A2(\gpout0.hpos[3] ),
    .B1(\gpout0.hpos[2] ),
    .B2(_04041_),
    .C1(_04059_),
    .X(_04060_));
 sky130_fd_sc_hd__a221o_1 _11342_ (.A1(_04055_),
    .A2(\gpout0.hpos[3] ),
    .B1(\gpout0.hpos[4] ),
    .B2(_04054_),
    .C1(_04060_),
    .X(_04061_));
 sky130_fd_sc_hd__o221a_1 _11343_ (.A1(_04053_),
    .A2(_03780_),
    .B1(\gpout0.hpos[4] ),
    .B2(_04054_),
    .C1(_04061_),
    .X(_04062_));
 sky130_fd_sc_hd__a221o_1 _11344_ (.A1(\rbzero.row_render.size[6] ),
    .A2(_03783_),
    .B1(_03780_),
    .B2(_04053_),
    .C1(_04062_),
    .X(_04063_));
 sky130_fd_sc_hd__o221a_1 _11345_ (.A1(\rbzero.row_render.size[6] ),
    .A2(_03783_),
    .B1(_03290_),
    .B2(_04052_),
    .C1(_04063_),
    .X(_04064_));
 sky130_fd_sc_hd__and2_1 _11346_ (.A(_03290_),
    .B(_04052_),
    .X(_04065_));
 sky130_fd_sc_hd__o22a_1 _11347_ (.A1(_03293_),
    .A2(_04050_),
    .B1(_04064_),
    .B2(_04065_),
    .X(_04066_));
 sky130_fd_sc_hd__a221o_1 _11348_ (.A1(_03293_),
    .A2(_04050_),
    .B1(_04051_),
    .B2(\gpout0.hpos[9] ),
    .C1(_04066_),
    .X(_04067_));
 sky130_fd_sc_hd__nand2_1 _11349_ (.A(\rbzero.row_render.size[9] ),
    .B(_04048_),
    .Y(_04068_));
 sky130_fd_sc_hd__o21a_1 _11350_ (.A1(_03295_),
    .A2(_04051_),
    .B1(_04068_),
    .X(_04069_));
 sky130_fd_sc_hd__nor3_1 _11351_ (.A(\rbzero.row_render.size[8] ),
    .B(\rbzero.row_render.size[7] ),
    .C(_04046_),
    .Y(_04070_));
 sky130_fd_sc_hd__nor2_1 _11352_ (.A(_04047_),
    .B(_04070_),
    .Y(_04071_));
 sky130_fd_sc_hd__xnor2_1 _11353_ (.A(\rbzero.row_render.size[7] ),
    .B(_04046_),
    .Y(_04072_));
 sky130_fd_sc_hd__a22o_1 _11354_ (.A1(_03290_),
    .A2(_04072_),
    .B1(_04071_),
    .B2(_03293_),
    .X(_04073_));
 sky130_fd_sc_hd__nor2_1 _11355_ (.A(\rbzero.row_render.size[6] ),
    .B(_04045_),
    .Y(_04074_));
 sky130_fd_sc_hd__nor2_1 _11356_ (.A(_04046_),
    .B(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__o21ai_1 _11357_ (.A1(\rbzero.row_render.size[4] ),
    .A2(_04044_),
    .B1(\rbzero.row_render.size[5] ),
    .Y(_04076_));
 sky130_fd_sc_hd__nand2_1 _11358_ (.A(_04045_),
    .B(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hd__clkbuf_4 _11359_ (.A(\gpout0.hpos[4] ),
    .X(_04078_));
 sky130_fd_sc_hd__xnor2_1 _11360_ (.A(\rbzero.row_render.size[4] ),
    .B(_04044_),
    .Y(_04079_));
 sky130_fd_sc_hd__clkbuf_4 _11361_ (.A(\gpout0.hpos[3] ),
    .X(_04080_));
 sky130_fd_sc_hd__nand2_1 _11362_ (.A(\rbzero.row_render.size[3] ),
    .B(_04043_),
    .Y(_04081_));
 sky130_fd_sc_hd__nand2_1 _11363_ (.A(_04044_),
    .B(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__or2_1 _11364_ (.A(_04041_),
    .B(_04042_),
    .X(_04083_));
 sky130_fd_sc_hd__nand2_1 _11365_ (.A(_04043_),
    .B(_04083_),
    .Y(_04084_));
 sky130_fd_sc_hd__and2_1 _11366_ (.A(\gpout0.hpos[1] ),
    .B(\gpout0.hpos[0] ),
    .X(_04085_));
 sky130_fd_sc_hd__or2_1 _11367_ (.A(\rbzero.row_render.size[0] ),
    .B(\gpout0.hpos[1] ),
    .X(_04086_));
 sky130_fd_sc_hd__or2_1 _11368_ (.A(\gpout0.hpos[1] ),
    .B(\gpout0.hpos[0] ),
    .X(_04087_));
 sky130_fd_sc_hd__a31o_1 _11369_ (.A1(\rbzero.row_render.size[1] ),
    .A2(_04086_),
    .A3(_04087_),
    .B1(_04042_),
    .X(_04088_));
 sky130_fd_sc_hd__a211o_1 _11370_ (.A1(\rbzero.row_render.size[2] ),
    .A2(\gpout0.hpos[2] ),
    .B1(_04085_),
    .C1(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__o221a_1 _11371_ (.A1(\gpout0.hpos[3] ),
    .A2(_04082_),
    .B1(_04084_),
    .B2(\gpout0.hpos[2] ),
    .C1(_04089_),
    .X(_04090_));
 sky130_fd_sc_hd__a221o_1 _11372_ (.A1(_04080_),
    .A2(_04082_),
    .B1(_04079_),
    .B2(\gpout0.hpos[4] ),
    .C1(_04090_),
    .X(_04091_));
 sky130_fd_sc_hd__o221a_1 _11373_ (.A1(_04078_),
    .A2(_04079_),
    .B1(_04077_),
    .B2(_03780_),
    .C1(_04091_),
    .X(_04092_));
 sky130_fd_sc_hd__a221o_1 _11374_ (.A1(_03781_),
    .A2(_04077_),
    .B1(_04075_),
    .B2(_03783_),
    .C1(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__o221a_1 _11375_ (.A1(_03784_),
    .A2(_04075_),
    .B1(_04072_),
    .B2(_03290_),
    .C1(_04093_),
    .X(_04094_));
 sky130_fd_sc_hd__o22a_1 _11376_ (.A1(_03293_),
    .A2(_04071_),
    .B1(_04073_),
    .B2(_04094_),
    .X(_04095_));
 sky130_fd_sc_hd__o2bb2a_1 _11377_ (.A1_N(_04067_),
    .A2_N(_04069_),
    .B1(_04095_),
    .B2(_03295_),
    .X(_04096_));
 sky130_fd_sc_hd__or4_2 _11378_ (.A(\rbzero.row_render.size[10] ),
    .B(\rbzero.row_render.size[9] ),
    .C(_04047_),
    .D(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__a21oi_1 _11379_ (.A1(_04040_),
    .A2(_04097_),
    .B1(\rbzero.row_render.vinf ),
    .Y(_04098_));
 sky130_fd_sc_hd__a221o_4 _11380_ (.A1(\rbzero.floor_leak[5] ),
    .A2(_03896_),
    .B1(_04036_),
    .B2(_04037_),
    .C1(_04098_),
    .X(_04099_));
 sky130_fd_sc_hd__mux2_1 _11381_ (.A0(_04028_),
    .A1(_04031_),
    .S(_04099_),
    .X(_04100_));
 sky130_fd_sc_hd__clkbuf_4 _11382_ (.A(\gpout0.vpos[3] ),
    .X(_04101_));
 sky130_fd_sc_hd__inv_2 _11383_ (.A(\gpout0.vpos[4] ),
    .Y(_04102_));
 sky130_fd_sc_hd__or2_2 _11384_ (.A(\gpout0.vpos[5] ),
    .B(_04102_),
    .X(_04103_));
 sky130_fd_sc_hd__buf_2 _11385_ (.A(\gpout0.vpos[5] ),
    .X(_04104_));
 sky130_fd_sc_hd__nand2_1 _11386_ (.A(_04104_),
    .B(_04101_),
    .Y(_04105_));
 sky130_fd_sc_hd__clkbuf_4 _11387_ (.A(\gpout0.vpos[4] ),
    .X(_04106_));
 sky130_fd_sc_hd__nand2_1 _11388_ (.A(\gpout0.hpos[2] ),
    .B(_04085_),
    .Y(_04107_));
 sky130_fd_sc_hd__o31a_2 _11389_ (.A1(\gpout0.vpos[2] ),
    .A2(\gpout0.vpos[1] ),
    .A3(\gpout0.vpos[0] ),
    .B1(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__o221ai_4 _11390_ (.A1(_04101_),
    .A2(_04103_),
    .B1(_04105_),
    .B2(_04106_),
    .C1(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__buf_2 _11391_ (.A(\gpout0.vpos[9] ),
    .X(_04110_));
 sky130_fd_sc_hd__clkinv_2 _11392_ (.A(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__and3_1 _11393_ (.A(\gpout0.vpos[8] ),
    .B(\gpout0.vpos[7] ),
    .C(\gpout0.vpos[6] ),
    .X(_04112_));
 sky130_fd_sc_hd__clkbuf_2 _11394_ (.A(_04112_),
    .X(_04113_));
 sky130_fd_sc_hd__nand2_1 _11395_ (.A(_04104_),
    .B(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hd__nand2_4 _11396_ (.A(_04111_),
    .B(_04114_),
    .Y(_04115_));
 sky130_fd_sc_hd__o21a_2 _11397_ (.A1(_03291_),
    .A2(_03294_),
    .B1(_03295_),
    .X(_04116_));
 sky130_fd_sc_hd__a211o_1 _11398_ (.A1(_03826_),
    .A2(_04109_),
    .B1(_04115_),
    .C1(_04116_),
    .X(_04117_));
 sky130_fd_sc_hd__o21bai_4 _11399_ (.A1(_03826_),
    .A2(_04100_),
    .B1_N(_04117_),
    .Y(_04118_));
 sky130_fd_sc_hd__inv_2 _11400_ (.A(_04118_),
    .Y(o_rgb[6]));
 sky130_fd_sc_hd__clkbuf_4 _11401_ (.A(_03934_),
    .X(_04119_));
 sky130_fd_sc_hd__mux2_1 _11402_ (.A0(\rbzero.tex_r1[49] ),
    .A1(\rbzero.tex_r1[48] ),
    .S(_04119_),
    .X(_04120_));
 sky130_fd_sc_hd__mux2_1 _11403_ (.A0(\rbzero.tex_r1[51] ),
    .A1(\rbzero.tex_r1[50] ),
    .S(_04119_),
    .X(_04121_));
 sky130_fd_sc_hd__mux2_1 _11404_ (.A0(_04120_),
    .A1(_04121_),
    .S(_03909_),
    .X(_04122_));
 sky130_fd_sc_hd__mux2_1 _11405_ (.A0(\rbzero.tex_r1[55] ),
    .A1(\rbzero.tex_r1[54] ),
    .S(_04119_),
    .X(_04123_));
 sky130_fd_sc_hd__mux2_1 _11406_ (.A0(\rbzero.tex_r1[53] ),
    .A1(\rbzero.tex_r1[52] ),
    .S(_04119_),
    .X(_04124_));
 sky130_fd_sc_hd__mux2_1 _11407_ (.A0(_04123_),
    .A1(_04124_),
    .S(_03942_),
    .X(_04125_));
 sky130_fd_sc_hd__mux2_1 _11408_ (.A0(_04122_),
    .A1(_04125_),
    .S(_03923_),
    .X(_04126_));
 sky130_fd_sc_hd__mux2_1 _11409_ (.A0(\rbzero.tex_r1[63] ),
    .A1(\rbzero.tex_r1[62] ),
    .S(_03935_),
    .X(_04127_));
 sky130_fd_sc_hd__mux2_1 _11410_ (.A0(\rbzero.tex_r1[61] ),
    .A1(\rbzero.tex_r1[60] ),
    .S(_03935_),
    .X(_04128_));
 sky130_fd_sc_hd__mux2_1 _11411_ (.A0(_04127_),
    .A1(_04128_),
    .S(_03942_),
    .X(_04129_));
 sky130_fd_sc_hd__mux2_1 _11412_ (.A0(\rbzero.tex_r1[57] ),
    .A1(\rbzero.tex_r1[56] ),
    .S(_03935_),
    .X(_04130_));
 sky130_fd_sc_hd__and2_1 _11413_ (.A(\rbzero.tex_r1[58] ),
    .B(_03925_),
    .X(_04131_));
 sky130_fd_sc_hd__a31o_1 _11414_ (.A1(\rbzero.tex_r1[59] ),
    .A2(_03938_),
    .A3(_03940_),
    .B1(_03915_),
    .X(_04132_));
 sky130_fd_sc_hd__o221a_1 _11415_ (.A1(_03910_),
    .A2(_04130_),
    .B1(_04131_),
    .B2(_04132_),
    .C1(_03945_),
    .X(_04133_));
 sky130_fd_sc_hd__a211o_1 _11416_ (.A1(_03921_),
    .A2(_04129_),
    .B1(_04133_),
    .C1(_03950_),
    .X(_04134_));
 sky130_fd_sc_hd__o211a_1 _11417_ (.A1(_03899_),
    .A2(_04126_),
    .B1(_04134_),
    .C1(_03954_),
    .X(_04135_));
 sky130_fd_sc_hd__mux2_1 _11418_ (.A0(\rbzero.tex_r1[45] ),
    .A1(\rbzero.tex_r1[44] ),
    .S(_03936_),
    .X(_04136_));
 sky130_fd_sc_hd__and2_1 _11419_ (.A(\rbzero.tex_r1[46] ),
    .B(_04013_),
    .X(_04137_));
 sky130_fd_sc_hd__a31o_1 _11420_ (.A1(\rbzero.tex_r1[47] ),
    .A2(_03939_),
    .A3(_03941_),
    .B1(_04014_),
    .X(_04138_));
 sky130_fd_sc_hd__o221a_1 _11421_ (.A1(_03932_),
    .A2(_04136_),
    .B1(_04137_),
    .B2(_04138_),
    .C1(_03923_),
    .X(_04139_));
 sky130_fd_sc_hd__mux2_1 _11422_ (.A0(\rbzero.tex_r1[43] ),
    .A1(\rbzero.tex_r1[42] ),
    .S(_03980_),
    .X(_04140_));
 sky130_fd_sc_hd__and2_1 _11423_ (.A(\rbzero.tex_r1[40] ),
    .B(_03959_),
    .X(_04141_));
 sky130_fd_sc_hd__clkbuf_4 _11424_ (.A(_03938_),
    .X(_04142_));
 sky130_fd_sc_hd__buf_2 _11425_ (.A(_04142_),
    .X(_04143_));
 sky130_fd_sc_hd__clkbuf_4 _11426_ (.A(_03940_),
    .X(_04144_));
 sky130_fd_sc_hd__buf_2 _11427_ (.A(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__a31o_1 _11428_ (.A1(\rbzero.tex_r1[41] ),
    .A2(_04143_),
    .A3(_04145_),
    .B1(_03910_),
    .X(_04146_));
 sky130_fd_sc_hd__o221a_1 _11429_ (.A1(_03968_),
    .A2(_04140_),
    .B1(_04141_),
    .B2(_04146_),
    .C1(_03972_),
    .X(_04147_));
 sky130_fd_sc_hd__buf_4 _11430_ (.A(_03934_),
    .X(_04148_));
 sky130_fd_sc_hd__mux2_1 _11431_ (.A0(\rbzero.tex_r1[39] ),
    .A1(\rbzero.tex_r1[38] ),
    .S(_04148_),
    .X(_04149_));
 sky130_fd_sc_hd__mux2_1 _11432_ (.A0(\rbzero.tex_r1[37] ),
    .A1(\rbzero.tex_r1[36] ),
    .S(_04148_),
    .X(_04150_));
 sky130_fd_sc_hd__mux2_1 _11433_ (.A0(_04149_),
    .A1(_04150_),
    .S(_04014_),
    .X(_04151_));
 sky130_fd_sc_hd__mux2_1 _11434_ (.A0(\rbzero.tex_r1[33] ),
    .A1(\rbzero.tex_r1[32] ),
    .S(_04148_),
    .X(_04152_));
 sky130_fd_sc_hd__and3_1 _11435_ (.A(\rbzero.tex_r1[35] ),
    .B(_03938_),
    .C(_03940_),
    .X(_04153_));
 sky130_fd_sc_hd__a21o_1 _11436_ (.A1(\rbzero.tex_r1[34] ),
    .A2(_03925_),
    .B1(_03915_),
    .X(_04154_));
 sky130_fd_sc_hd__o221a_1 _11437_ (.A1(_03910_),
    .A2(_04152_),
    .B1(_04153_),
    .B2(_04154_),
    .C1(_03945_),
    .X(_04155_));
 sky130_fd_sc_hd__a211o_1 _11438_ (.A1(_03921_),
    .A2(_04151_),
    .B1(_04155_),
    .C1(_03898_),
    .X(_04156_));
 sky130_fd_sc_hd__o311a_1 _11439_ (.A1(_03956_),
    .A2(_04139_),
    .A3(_04147_),
    .B1(_04156_),
    .C1(_03985_),
    .X(_04157_));
 sky130_fd_sc_hd__mux2_1 _11440_ (.A0(\rbzero.tex_r1[19] ),
    .A1(\rbzero.tex_r1[18] ),
    .S(_04000_),
    .X(_04158_));
 sky130_fd_sc_hd__mux2_1 _11441_ (.A0(\rbzero.tex_r1[17] ),
    .A1(\rbzero.tex_r1[16] ),
    .S(_04148_),
    .X(_04159_));
 sky130_fd_sc_hd__mux2_1 _11442_ (.A0(_04158_),
    .A1(_04159_),
    .S(_04014_),
    .X(_04160_));
 sky130_fd_sc_hd__mux2_1 _11443_ (.A0(\rbzero.tex_r1[21] ),
    .A1(\rbzero.tex_r1[20] ),
    .S(_04000_),
    .X(_04161_));
 sky130_fd_sc_hd__mux2_1 _11444_ (.A0(\rbzero.tex_r1[23] ),
    .A1(\rbzero.tex_r1[22] ),
    .S(_04148_),
    .X(_04162_));
 sky130_fd_sc_hd__mux2_1 _11445_ (.A0(_04161_),
    .A1(_04162_),
    .S(_03910_),
    .X(_04163_));
 sky130_fd_sc_hd__mux2_1 _11446_ (.A0(_04160_),
    .A1(_04163_),
    .S(_03923_),
    .X(_04164_));
 sky130_fd_sc_hd__mux2_1 _11447_ (.A0(\rbzero.tex_r1[27] ),
    .A1(\rbzero.tex_r1[26] ),
    .S(_03904_),
    .X(_04165_));
 sky130_fd_sc_hd__mux2_1 _11448_ (.A0(\rbzero.tex_r1[25] ),
    .A1(\rbzero.tex_r1[24] ),
    .S(_03904_),
    .X(_04166_));
 sky130_fd_sc_hd__mux2_1 _11449_ (.A0(_04165_),
    .A1(_04166_),
    .S(_03916_),
    .X(_04167_));
 sky130_fd_sc_hd__buf_4 _11450_ (.A(_03903_),
    .X(_04168_));
 sky130_fd_sc_hd__mux2_1 _11451_ (.A0(\rbzero.tex_r1[29] ),
    .A1(\rbzero.tex_r1[28] ),
    .S(_04168_),
    .X(_04169_));
 sky130_fd_sc_hd__and2_1 _11452_ (.A(\rbzero.tex_r1[30] ),
    .B(_03961_),
    .X(_04170_));
 sky130_fd_sc_hd__a31o_1 _11453_ (.A1(\rbzero.tex_r1[31] ),
    .A2(_04142_),
    .A3(_04144_),
    .B1(_03929_),
    .X(_04171_));
 sky130_fd_sc_hd__o221a_1 _11454_ (.A1(_03957_),
    .A2(_04169_),
    .B1(_04170_),
    .B2(_04171_),
    .C1(_03923_),
    .X(_04172_));
 sky130_fd_sc_hd__a211o_1 _11455_ (.A1(_03972_),
    .A2(_04167_),
    .B1(_04172_),
    .C1(_03950_),
    .X(_04173_));
 sky130_fd_sc_hd__o211a_1 _11456_ (.A1(_03900_),
    .A2(_04164_),
    .B1(_04173_),
    .C1(_03954_),
    .X(_04174_));
 sky130_fd_sc_hd__mux2_1 _11457_ (.A0(\rbzero.tex_r1[15] ),
    .A1(\rbzero.tex_r1[14] ),
    .S(_04168_),
    .X(_04175_));
 sky130_fd_sc_hd__mux2_1 _11458_ (.A0(\rbzero.tex_r1[13] ),
    .A1(\rbzero.tex_r1[12] ),
    .S(_04168_),
    .X(_04176_));
 sky130_fd_sc_hd__mux2_1 _11459_ (.A0(_04175_),
    .A1(_04176_),
    .S(_03916_),
    .X(_04177_));
 sky130_fd_sc_hd__mux2_1 _11460_ (.A0(\rbzero.tex_r1[9] ),
    .A1(\rbzero.tex_r1[8] ),
    .S(_04168_),
    .X(_04178_));
 sky130_fd_sc_hd__and3_1 _11461_ (.A(\rbzero.tex_r1[11] ),
    .B(_04142_),
    .C(_04144_),
    .X(_04179_));
 sky130_fd_sc_hd__a21o_1 _11462_ (.A1(\rbzero.tex_r1[10] ),
    .A2(_03961_),
    .B1(_03929_),
    .X(_04180_));
 sky130_fd_sc_hd__o221a_1 _11463_ (.A1(_03957_),
    .A2(_04178_),
    .B1(_04179_),
    .B2(_04180_),
    .C1(_03946_),
    .X(_04181_));
 sky130_fd_sc_hd__a211o_1 _11464_ (.A1(_03924_),
    .A2(_04177_),
    .B1(_04181_),
    .C1(_03950_),
    .X(_04182_));
 sky130_fd_sc_hd__mux2_1 _11465_ (.A0(\rbzero.tex_r1[5] ),
    .A1(\rbzero.tex_r1[4] ),
    .S(_04168_),
    .X(_04183_));
 sky130_fd_sc_hd__mux2_1 _11466_ (.A0(\rbzero.tex_r1[7] ),
    .A1(\rbzero.tex_r1[6] ),
    .S(_04168_),
    .X(_04184_));
 sky130_fd_sc_hd__mux2_1 _11467_ (.A0(_04183_),
    .A1(_04184_),
    .S(_03910_),
    .X(_04185_));
 sky130_fd_sc_hd__and3_1 _11468_ (.A(\rbzero.tex_r1[3] ),
    .B(_04142_),
    .C(_04144_),
    .X(_04186_));
 sky130_fd_sc_hd__a21o_1 _11469_ (.A1(\rbzero.tex_r1[2] ),
    .A2(_03961_),
    .B1(_03929_),
    .X(_04187_));
 sky130_fd_sc_hd__mux2_1 _11470_ (.A0(\rbzero.tex_r1[1] ),
    .A1(\rbzero.tex_r1[0] ),
    .S(_04168_),
    .X(_04188_));
 sky130_fd_sc_hd__o221a_1 _11471_ (.A1(_04186_),
    .A2(_04187_),
    .B1(_04188_),
    .B2(_03957_),
    .C1(_03946_),
    .X(_04189_));
 sky130_fd_sc_hd__a211o_1 _11472_ (.A1(_03924_),
    .A2(_04185_),
    .B1(_04189_),
    .C1(_03899_),
    .X(_04190_));
 sky130_fd_sc_hd__a31o_1 _11473_ (.A1(_03985_),
    .A2(_04182_),
    .A3(_04190_),
    .B1(_04026_),
    .X(_04191_));
 sky130_fd_sc_hd__o32a_1 _11474_ (.A1(_03896_),
    .A2(_04135_),
    .A3(_04157_),
    .B1(_04174_),
    .B2(_04191_),
    .X(_04192_));
 sky130_fd_sc_hd__mux2_1 _11475_ (.A0(\rbzero.color_sky[1] ),
    .A1(\rbzero.color_floor[1] ),
    .S(_04030_),
    .X(_04193_));
 sky130_fd_sc_hd__mux2_1 _11476_ (.A0(_04192_),
    .A1(_04193_),
    .S(_04099_),
    .X(_04194_));
 sky130_fd_sc_hd__a21oi_1 _11477_ (.A1(\gpout0.hpos[3] ),
    .A2(_03804_),
    .B1(\gpout0.hpos[4] ),
    .Y(_04195_));
 sky130_fd_sc_hd__or2_1 _11478_ (.A(_03806_),
    .B(_04195_),
    .X(_04196_));
 sky130_fd_sc_hd__nand2_1 _11479_ (.A(_03802_),
    .B(_03824_),
    .Y(_04197_));
 sky130_fd_sc_hd__xnor2_1 _11480_ (.A(\gpout0.hpos[3] ),
    .B(_03804_),
    .Y(_04198_));
 sky130_fd_sc_hd__or2b_1 _11481_ (.A(_04197_),
    .B_N(_04198_),
    .X(_04199_));
 sky130_fd_sc_hd__nor2_1 _11482_ (.A(_04196_),
    .B(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__nand2_1 _11483_ (.A(_03780_),
    .B(_04200_),
    .Y(_04201_));
 sky130_fd_sc_hd__nand3_1 _11484_ (.A(_03783_),
    .B(\gpout0.hpos[5] ),
    .C(_03806_),
    .Y(_04202_));
 sky130_fd_sc_hd__nand2_2 _11485_ (.A(_03823_),
    .B(_04202_),
    .Y(_04203_));
 sky130_fd_sc_hd__nand2_1 _11486_ (.A(_03788_),
    .B(_04202_),
    .Y(_04204_));
 sky130_fd_sc_hd__nor2_1 _11487_ (.A(_03788_),
    .B(_04202_),
    .Y(_04205_));
 sky130_fd_sc_hd__nand2_2 _11488_ (.A(_03293_),
    .B(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hd__o21ai_4 _11489_ (.A1(_03293_),
    .A2(_04204_),
    .B1(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hd__nand2_2 _11490_ (.A(_04203_),
    .B(_04207_),
    .Y(_04208_));
 sky130_fd_sc_hd__nor2_2 _11491_ (.A(_04201_),
    .B(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__xor2_1 _11492_ (.A(\gpout0.hpos[5] ),
    .B(_03806_),
    .X(_04210_));
 sky130_fd_sc_hd__a21boi_1 _11493_ (.A1(_03290_),
    .A2(_03823_),
    .B1_N(_04204_),
    .Y(_04211_));
 sky130_fd_sc_hd__or4b_1 _11494_ (.A(_04199_),
    .B(_04210_),
    .C(_04211_),
    .D_N(_04196_),
    .X(_04212_));
 sky130_fd_sc_hd__nor2_1 _11495_ (.A(_04203_),
    .B(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__and2_2 _11496_ (.A(_04213_),
    .B(_04207_),
    .X(_04214_));
 sky130_fd_sc_hd__or2_1 _11497_ (.A(_04198_),
    .B(_04197_),
    .X(_04215_));
 sky130_fd_sc_hd__or3b_1 _11498_ (.A(_04210_),
    .B(_04215_),
    .C_N(\gpout0.hpos[4] ),
    .X(_04216_));
 sky130_fd_sc_hd__nor2_1 _11499_ (.A(_04203_),
    .B(_04216_),
    .Y(_04217_));
 sky130_fd_sc_hd__and2_2 _11500_ (.A(_04217_),
    .B(_04207_),
    .X(_04218_));
 sky130_fd_sc_hd__a22o_1 _11501_ (.A1(\rbzero.debug_overlay.facingX[-5] ),
    .A2(_04214_),
    .B1(_04218_),
    .B2(\rbzero.debug_overlay.facingX[-8] ),
    .X(_04219_));
 sky130_fd_sc_hd__xnor2_1 _11502_ (.A(_03780_),
    .B(_03806_),
    .Y(_04220_));
 sky130_fd_sc_hd__nor2_1 _11503_ (.A(_04215_),
    .B(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__a211o_1 _11504_ (.A1(_03803_),
    .A2(_04200_),
    .B1(_04217_),
    .C1(_04221_),
    .X(_04222_));
 sky130_fd_sc_hd__nor3_1 _11505_ (.A(_03780_),
    .B(\gpout0.hpos[4] ),
    .C(_04215_),
    .Y(_04223_));
 sky130_fd_sc_hd__inv_2 _11506_ (.A(_03783_),
    .Y(_04224_));
 sky130_fd_sc_hd__or3b_2 _11507_ (.A(_04199_),
    .B(_04220_),
    .C_N(_04196_),
    .X(_04225_));
 sky130_fd_sc_hd__nor2_1 _11508_ (.A(_04224_),
    .B(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__a211o_1 _11509_ (.A1(_03783_),
    .A2(_04223_),
    .B1(_04213_),
    .C1(_04226_),
    .X(_04227_));
 sky130_fd_sc_hd__and2b_1 _11510_ (.A_N(_04205_),
    .B(_04204_),
    .X(_04228_));
 sky130_fd_sc_hd__nand2_1 _11511_ (.A(_03293_),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__o21ba_1 _11512_ (.A1(_04222_),
    .A2(_04227_),
    .B1_N(_04229_),
    .X(_04230_));
 sky130_fd_sc_hd__nor2_1 _11513_ (.A(_04212_),
    .B(_04208_),
    .Y(_04231_));
 sky130_fd_sc_hd__and2b_1 _11514_ (.A_N(_03780_),
    .B(_04200_),
    .X(_04232_));
 sky130_fd_sc_hd__and2_1 _11515_ (.A(_04203_),
    .B(_04207_),
    .X(_04233_));
 sky130_fd_sc_hd__and2_1 _11516_ (.A(_04232_),
    .B(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__and2_1 _11517_ (.A(_04223_),
    .B(_04233_),
    .X(_04235_));
 sky130_fd_sc_hd__or4_2 _11518_ (.A(_04230_),
    .B(_04231_),
    .C(_04234_),
    .D(_04235_),
    .X(_04236_));
 sky130_fd_sc_hd__and3_2 _11519_ (.A(_03783_),
    .B(_04223_),
    .C(_04207_),
    .X(_04237_));
 sky130_fd_sc_hd__and3_2 _11520_ (.A(_03783_),
    .B(_04232_),
    .C(_04207_),
    .X(_04238_));
 sky130_fd_sc_hd__a22o_1 _11521_ (.A1(\rbzero.debug_overlay.facingX[-6] ),
    .A2(_04237_),
    .B1(_04238_),
    .B2(\rbzero.debug_overlay.facingX[-7] ),
    .X(_04239_));
 sky130_fd_sc_hd__and2_2 _11522_ (.A(_04226_),
    .B(_04207_),
    .X(_04240_));
 sky130_fd_sc_hd__nand2_1 _11523_ (.A(_04078_),
    .B(_04221_),
    .Y(_04241_));
 sky130_fd_sc_hd__nor2_2 _11524_ (.A(_04208_),
    .B(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__nor2_2 _11525_ (.A(_04216_),
    .B(_04208_),
    .Y(_04243_));
 sky130_fd_sc_hd__nor2_4 _11526_ (.A(_04225_),
    .B(_04208_),
    .Y(_04244_));
 sky130_fd_sc_hd__and4bb_2 _11527_ (.A_N(\gpout0.hpos[4] ),
    .B_N(_04215_),
    .C(_04233_),
    .D(_03780_),
    .X(_04245_));
 sky130_fd_sc_hd__inv_2 _11528_ (.A(\gpout0.vpos[3] ),
    .Y(_04246_));
 sky130_fd_sc_hd__a211o_1 _11529_ (.A1(\rbzero.debug_overlay.facingX[-2] ),
    .A2(_04245_),
    .B1(_04103_),
    .C1(_04246_),
    .X(_04247_));
 sky130_fd_sc_hd__a221o_1 _11530_ (.A1(\rbzero.debug_overlay.facingX[0] ),
    .A2(_04243_),
    .B1(_04244_),
    .B2(\rbzero.debug_overlay.facingX[-1] ),
    .C1(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__a221o_1 _11531_ (.A1(\rbzero.debug_overlay.facingX[-9] ),
    .A2(_04240_),
    .B1(_04242_),
    .B2(\rbzero.debug_overlay.facingX[-4] ),
    .C1(_04248_),
    .X(_04249_));
 sky130_fd_sc_hd__a211o_1 _11532_ (.A1(\rbzero.debug_overlay.facingX[10] ),
    .A2(_04236_),
    .B1(_04239_),
    .C1(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__a211o_1 _11533_ (.A1(\rbzero.debug_overlay.facingX[-3] ),
    .A2(_04209_),
    .B1(_04219_),
    .C1(_04250_),
    .X(_04251_));
 sky130_fd_sc_hd__nor2_2 _11534_ (.A(_04104_),
    .B(_04102_),
    .Y(_04252_));
 sky130_fd_sc_hd__a22o_1 _11535_ (.A1(\rbzero.debug_overlay.vplaneX[-5] ),
    .A2(_04214_),
    .B1(_04237_),
    .B2(\rbzero.debug_overlay.vplaneX[-6] ),
    .X(_04253_));
 sky130_fd_sc_hd__a22o_1 _11536_ (.A1(\rbzero.debug_overlay.vplaneX[-4] ),
    .A2(_04242_),
    .B1(_04209_),
    .B2(\rbzero.debug_overlay.vplaneX[-3] ),
    .X(_04254_));
 sky130_fd_sc_hd__a221o_1 _11537_ (.A1(\rbzero.debug_overlay.vplaneX[-2] ),
    .A2(_04245_),
    .B1(_04243_),
    .B2(\rbzero.debug_overlay.vplaneX[0] ),
    .C1(\gpout0.vpos[3] ),
    .X(_04255_));
 sky130_fd_sc_hd__a221o_1 _11538_ (.A1(\rbzero.debug_overlay.vplaneX[-8] ),
    .A2(_04218_),
    .B1(_04244_),
    .B2(\rbzero.debug_overlay.vplaneX[-1] ),
    .C1(_04255_),
    .X(_04256_));
 sky130_fd_sc_hd__a211o_1 _11539_ (.A1(\rbzero.debug_overlay.vplaneX[-7] ),
    .A2(_04238_),
    .B1(_04254_),
    .C1(_04256_),
    .X(_04257_));
 sky130_fd_sc_hd__a211o_1 _11540_ (.A1(\rbzero.debug_overlay.vplaneX[-9] ),
    .A2(_04240_),
    .B1(_04253_),
    .C1(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__a21o_1 _11541_ (.A1(\rbzero.debug_overlay.vplaneX[10] ),
    .A2(_04236_),
    .B1(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__buf_2 _11542_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .X(_04260_));
 sky130_fd_sc_hd__a22o_1 _11543_ (.A1(\rbzero.debug_overlay.vplaneY[-4] ),
    .A2(_04242_),
    .B1(_04245_),
    .B2(_04260_),
    .X(_04261_));
 sky130_fd_sc_hd__a221o_1 _11544_ (.A1(\rbzero.debug_overlay.vplaneY[-3] ),
    .A2(_04209_),
    .B1(_04243_),
    .B2(\rbzero.debug_overlay.vplaneY[0] ),
    .C1(_04261_),
    .X(_04262_));
 sky130_fd_sc_hd__a221o_1 _11545_ (.A1(\rbzero.debug_overlay.vplaneY[-7] ),
    .A2(_04238_),
    .B1(_04244_),
    .B2(\rbzero.debug_overlay.vplaneY[-1] ),
    .C1(_04246_),
    .X(_04263_));
 sky130_fd_sc_hd__a22o_1 _11546_ (.A1(\rbzero.debug_overlay.vplaneY[-5] ),
    .A2(_04214_),
    .B1(_04237_),
    .B2(\rbzero.debug_overlay.vplaneY[-6] ),
    .X(_04264_));
 sky130_fd_sc_hd__a221o_1 _11547_ (.A1(\rbzero.debug_overlay.vplaneY[-9] ),
    .A2(_04240_),
    .B1(_04218_),
    .B2(\rbzero.debug_overlay.vplaneY[-8] ),
    .C1(_04264_),
    .X(_04265_));
 sky130_fd_sc_hd__a211o_1 _11548_ (.A1(\rbzero.debug_overlay.vplaneY[10] ),
    .A2(_04236_),
    .B1(_04263_),
    .C1(_04265_),
    .X(_04266_));
 sky130_fd_sc_hd__o211a_1 _11549_ (.A1(_04262_),
    .A2(_04266_),
    .B1(\gpout0.vpos[5] ),
    .C1(_04106_),
    .X(_04267_));
 sky130_fd_sc_hd__a22o_1 _11550_ (.A1(\rbzero.debug_overlay.facingY[-9] ),
    .A2(_04240_),
    .B1(_04218_),
    .B2(\rbzero.debug_overlay.facingY[-8] ),
    .X(_04268_));
 sky130_fd_sc_hd__a221o_1 _11551_ (.A1(\rbzero.debug_overlay.facingY[-4] ),
    .A2(_04242_),
    .B1(_04209_),
    .B2(\rbzero.debug_overlay.facingY[-3] ),
    .C1(_04268_),
    .X(_04269_));
 sky130_fd_sc_hd__a22o_1 _11552_ (.A1(\rbzero.debug_overlay.facingY[-2] ),
    .A2(_04245_),
    .B1(_04243_),
    .B2(\rbzero.debug_overlay.facingY[0] ),
    .X(_04270_));
 sky130_fd_sc_hd__a221o_1 _11553_ (.A1(\rbzero.debug_overlay.facingY[-5] ),
    .A2(_04214_),
    .B1(_04244_),
    .B2(\rbzero.debug_overlay.facingY[-1] ),
    .C1(_04270_),
    .X(_04271_));
 sky130_fd_sc_hd__a221o_1 _11554_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(_04237_),
    .B1(_04238_),
    .B2(\rbzero.debug_overlay.facingY[-7] ),
    .C1(_04271_),
    .X(_04272_));
 sky130_fd_sc_hd__a21o_1 _11555_ (.A1(\rbzero.debug_overlay.facingY[10] ),
    .A2(_04236_),
    .B1(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__o2111a_1 _11556_ (.A1(_04269_),
    .A2(_04273_),
    .B1(\gpout0.vpos[5] ),
    .C1(_04102_),
    .D1(_04246_),
    .X(_04274_));
 sky130_fd_sc_hd__a221o_1 _11557_ (.A1(\gpout0.vpos[3] ),
    .A2(_04252_),
    .B1(_04259_),
    .B2(_04267_),
    .C1(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__a2bb2o_1 _11558_ (.A1_N(_04104_),
    .A2_N(_04106_),
    .B1(_04251_),
    .B2(_04275_),
    .X(_04276_));
 sky130_fd_sc_hd__a22o_1 _11559_ (.A1(\rbzero.debug_overlay.playerY[-5] ),
    .A2(_04214_),
    .B1(_04237_),
    .B2(\rbzero.debug_overlay.playerY[-6] ),
    .X(_04277_));
 sky130_fd_sc_hd__nor2_1 _11560_ (.A(_04229_),
    .B(_04241_),
    .Y(_04278_));
 sky130_fd_sc_hd__a22o_1 _11561_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_04231_),
    .B1(_04244_),
    .B2(\rbzero.debug_overlay.playerY[-1] ),
    .X(_04279_));
 sky130_fd_sc_hd__a221o_1 _11562_ (.A1(\rbzero.debug_overlay.playerY[-8] ),
    .A2(_04218_),
    .B1(_04278_),
    .B2(\rbzero.debug_overlay.playerY[4] ),
    .C1(_04279_),
    .X(_04280_));
 sky130_fd_sc_hd__a22o_1 _11563_ (.A1(\rbzero.debug_overlay.playerY[-4] ),
    .A2(_04242_),
    .B1(_04238_),
    .B2(\rbzero.debug_overlay.playerY[-7] ),
    .X(_04281_));
 sky130_fd_sc_hd__nor2_1 _11564_ (.A(_04229_),
    .B(_04201_),
    .Y(_04282_));
 sky130_fd_sc_hd__a22o_1 _11565_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_04235_),
    .B1(_04282_),
    .B2(\rbzero.debug_overlay.playerY[5] ),
    .X(_04283_));
 sky130_fd_sc_hd__or3_1 _11566_ (.A(\gpout0.vpos[5] ),
    .B(\gpout0.vpos[4] ),
    .C(_04246_),
    .X(_04284_));
 sky130_fd_sc_hd__a221o_1 _11567_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_04245_),
    .B1(_04243_),
    .B2(\rbzero.debug_overlay.playerY[0] ),
    .C1(_04284_),
    .X(_04285_));
 sky130_fd_sc_hd__a221o_1 _11568_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_04234_),
    .B1(_04209_),
    .B2(\rbzero.debug_overlay.playerY[-3] ),
    .C1(_04285_),
    .X(_04286_));
 sky130_fd_sc_hd__or4_1 _11569_ (.A(_04280_),
    .B(_04281_),
    .C(_04283_),
    .D(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__a211o_1 _11570_ (.A1(\rbzero.debug_overlay.playerY[-9] ),
    .A2(_04240_),
    .B1(_04277_),
    .C1(_04287_),
    .X(_04288_));
 sky130_fd_sc_hd__a22o_1 _11571_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_04214_),
    .B1(_04237_),
    .B2(\rbzero.debug_overlay.playerX[-6] ),
    .X(_04289_));
 sky130_fd_sc_hd__a22o_1 _11572_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_04235_),
    .B1(_04278_),
    .B2(\rbzero.debug_overlay.playerX[4] ),
    .X(_04290_));
 sky130_fd_sc_hd__a221o_1 _11573_ (.A1(\rbzero.debug_overlay.playerX[-4] ),
    .A2(_04242_),
    .B1(_04244_),
    .B2(\rbzero.debug_overlay.playerX[-1] ),
    .C1(_04290_),
    .X(_04291_));
 sky130_fd_sc_hd__a22o_1 _11574_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_04231_),
    .B1(_04209_),
    .B2(\rbzero.debug_overlay.playerX[-3] ),
    .X(_04292_));
 sky130_fd_sc_hd__a221o_1 _11575_ (.A1(\rbzero.debug_overlay.playerX[-8] ),
    .A2(_04218_),
    .B1(_04238_),
    .B2(\rbzero.debug_overlay.playerX[-7] ),
    .C1(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__a221o_1 _11576_ (.A1(\rbzero.debug_overlay.playerX[-2] ),
    .A2(_04245_),
    .B1(_04243_),
    .B2(\rbzero.debug_overlay.playerX[0] ),
    .C1(_03821_),
    .X(_04294_));
 sky130_fd_sc_hd__a221o_1 _11577_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_04234_),
    .B1(_04282_),
    .B2(\rbzero.debug_overlay.playerX[5] ),
    .C1(_04294_),
    .X(_04295_));
 sky130_fd_sc_hd__or3_1 _11578_ (.A(_04291_),
    .B(_04293_),
    .C(_04295_),
    .X(_04296_));
 sky130_fd_sc_hd__a211o_1 _11579_ (.A1(\rbzero.debug_overlay.playerX[-9] ),
    .A2(_04240_),
    .B1(_04289_),
    .C1(_04296_),
    .X(_04297_));
 sky130_fd_sc_hd__and3_1 _11580_ (.A(_04108_),
    .B(_04288_),
    .C(_04297_),
    .X(_04298_));
 sky130_fd_sc_hd__nand2_1 _11581_ (.A(_04276_),
    .B(_04298_),
    .Y(_04299_));
 sky130_fd_sc_hd__o311a_1 _11582_ (.A1(_03293_),
    .A2(_03296_),
    .A3(_03807_),
    .B1(_03826_),
    .C1(_04299_),
    .X(_04300_));
 sky130_fd_sc_hd__or3_1 _11583_ (.A(_04116_),
    .B(_04115_),
    .C(_04300_),
    .X(_04301_));
 sky130_fd_sc_hd__o21ba_1 _11584_ (.A1(_03826_),
    .A2(_04194_),
    .B1_N(_04301_),
    .X(_04302_));
 sky130_fd_sc_hd__buf_4 _11585_ (.A(_04302_),
    .X(o_rgb[7]));
 sky130_fd_sc_hd__mux2_1 _11586_ (.A0(\rbzero.tex_g0[19] ),
    .A1(\rbzero.tex_g0[18] ),
    .S(_04119_),
    .X(_04303_));
 sky130_fd_sc_hd__mux2_1 _11587_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_04119_),
    .X(_04304_));
 sky130_fd_sc_hd__mux2_1 _11588_ (.A0(_04303_),
    .A1(_04304_),
    .S(_03942_),
    .X(_04305_));
 sky130_fd_sc_hd__mux2_1 _11589_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(_04119_),
    .X(_04306_));
 sky130_fd_sc_hd__mux2_1 _11590_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(_04119_),
    .X(_04307_));
 sky130_fd_sc_hd__mux2_1 _11591_ (.A0(_04306_),
    .A1(_04307_),
    .S(_03909_),
    .X(_04308_));
 sky130_fd_sc_hd__mux2_1 _11592_ (.A0(_04305_),
    .A1(_04308_),
    .S(_03923_),
    .X(_04309_));
 sky130_fd_sc_hd__mux2_1 _11593_ (.A0(\rbzero.tex_g0[27] ),
    .A1(\rbzero.tex_g0[26] ),
    .S(_03935_),
    .X(_04310_));
 sky130_fd_sc_hd__mux2_1 _11594_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_03935_),
    .X(_04311_));
 sky130_fd_sc_hd__mux2_1 _11595_ (.A0(_04310_),
    .A1(_04311_),
    .S(_03942_),
    .X(_04312_));
 sky130_fd_sc_hd__mux2_1 _11596_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_03935_),
    .X(_04313_));
 sky130_fd_sc_hd__and2_1 _11597_ (.A(\rbzero.tex_g0[30] ),
    .B(_04168_),
    .X(_04314_));
 sky130_fd_sc_hd__a31o_1 _11598_ (.A1(\rbzero.tex_g0[31] ),
    .A2(_03938_),
    .A3(_03940_),
    .B1(_03915_),
    .X(_04315_));
 sky130_fd_sc_hd__o221a_1 _11599_ (.A1(_03910_),
    .A2(_04313_),
    .B1(_04314_),
    .B2(_04315_),
    .C1(_03920_),
    .X(_04316_));
 sky130_fd_sc_hd__a211o_1 _11600_ (.A1(_03972_),
    .A2(_04312_),
    .B1(_04316_),
    .C1(_03950_),
    .X(_04317_));
 sky130_fd_sc_hd__o211a_1 _11601_ (.A1(_03899_),
    .A2(_04309_),
    .B1(_04317_),
    .C1(_03954_),
    .X(_04318_));
 sky130_fd_sc_hd__and3_1 _11602_ (.A(\rbzero.tex_g0[3] ),
    .B(_03939_),
    .C(_03941_),
    .X(_04319_));
 sky130_fd_sc_hd__a21o_1 _11603_ (.A1(\rbzero.tex_g0[2] ),
    .A2(_04013_),
    .B1(_04014_),
    .X(_04320_));
 sky130_fd_sc_hd__mux2_1 _11604_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_03936_),
    .X(_04321_));
 sky130_fd_sc_hd__o221a_1 _11605_ (.A1(_04319_),
    .A2(_04320_),
    .B1(_04321_),
    .B2(_03932_),
    .C1(_03946_),
    .X(_04322_));
 sky130_fd_sc_hd__buf_4 _11606_ (.A(_03910_),
    .X(_04323_));
 sky130_fd_sc_hd__mux2_1 _11607_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_03936_),
    .X(_04324_));
 sky130_fd_sc_hd__and2_1 _11608_ (.A(\rbzero.tex_g0[6] ),
    .B(_04013_),
    .X(_04325_));
 sky130_fd_sc_hd__a31o_1 _11609_ (.A1(\rbzero.tex_g0[7] ),
    .A2(_03939_),
    .A3(_03941_),
    .B1(_04014_),
    .X(_04326_));
 sky130_fd_sc_hd__o221a_1 _11610_ (.A1(_04323_),
    .A2(_04324_),
    .B1(_04325_),
    .B2(_04326_),
    .C1(_03923_),
    .X(_04327_));
 sky130_fd_sc_hd__mux2_1 _11611_ (.A0(\rbzero.tex_g0[15] ),
    .A1(\rbzero.tex_g0[14] ),
    .S(_04148_),
    .X(_04328_));
 sky130_fd_sc_hd__mux2_1 _11612_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_04148_),
    .X(_04329_));
 sky130_fd_sc_hd__mux2_1 _11613_ (.A0(_04328_),
    .A1(_04329_),
    .S(_04014_),
    .X(_04330_));
 sky130_fd_sc_hd__mux2_1 _11614_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_04148_),
    .X(_04331_));
 sky130_fd_sc_hd__and3_1 _11615_ (.A(\rbzero.tex_g0[11] ),
    .B(_04142_),
    .C(_04144_),
    .X(_04332_));
 sky130_fd_sc_hd__a21o_1 _11616_ (.A1(\rbzero.tex_g0[10] ),
    .A2(_03974_),
    .B1(_03929_),
    .X(_04333_));
 sky130_fd_sc_hd__o221a_1 _11617_ (.A1(_03910_),
    .A2(_04331_),
    .B1(_04332_),
    .B2(_04333_),
    .C1(_03945_),
    .X(_04334_));
 sky130_fd_sc_hd__a211o_1 _11618_ (.A1(_03921_),
    .A2(_04330_),
    .B1(_04334_),
    .C1(_03950_),
    .X(_04335_));
 sky130_fd_sc_hd__o311a_1 _11619_ (.A1(_03899_),
    .A2(_04322_),
    .A3(_04327_),
    .B1(_03985_),
    .C1(_04335_),
    .X(_04336_));
 sky130_fd_sc_hd__mux2_1 _11620_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_04148_),
    .X(_04337_));
 sky130_fd_sc_hd__mux2_1 _11621_ (.A0(\rbzero.tex_g0[51] ),
    .A1(\rbzero.tex_g0[50] ),
    .S(_03935_),
    .X(_04338_));
 sky130_fd_sc_hd__mux2_1 _11622_ (.A0(_04337_),
    .A1(_04338_),
    .S(_03909_),
    .X(_04339_));
 sky130_fd_sc_hd__mux2_1 _11623_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(_04148_),
    .X(_04340_));
 sky130_fd_sc_hd__mux2_1 _11624_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(_03935_),
    .X(_04341_));
 sky130_fd_sc_hd__mux2_1 _11625_ (.A0(_04340_),
    .A1(_04341_),
    .S(_03942_),
    .X(_04342_));
 sky130_fd_sc_hd__mux2_1 _11626_ (.A0(_04339_),
    .A1(_04342_),
    .S(_03923_),
    .X(_04343_));
 sky130_fd_sc_hd__mux2_1 _11627_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(_04168_),
    .X(_04344_));
 sky130_fd_sc_hd__mux2_1 _11628_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_04168_),
    .X(_04345_));
 sky130_fd_sc_hd__mux2_1 _11629_ (.A0(_04344_),
    .A1(_04345_),
    .S(_04014_),
    .X(_04346_));
 sky130_fd_sc_hd__mux2_1 _11630_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(_04000_),
    .X(_04347_));
 sky130_fd_sc_hd__and2_1 _11631_ (.A(\rbzero.tex_g0[58] ),
    .B(_03974_),
    .X(_04348_));
 sky130_fd_sc_hd__a31o_1 _11632_ (.A1(\rbzero.tex_g0[59] ),
    .A2(_04142_),
    .A3(_04144_),
    .B1(_03929_),
    .X(_04349_));
 sky130_fd_sc_hd__o221a_1 _11633_ (.A1(_03957_),
    .A2(_04347_),
    .B1(_04348_),
    .B2(_04349_),
    .C1(_03945_),
    .X(_04350_));
 sky130_fd_sc_hd__a211o_1 _11634_ (.A1(_03921_),
    .A2(_04346_),
    .B1(_04350_),
    .C1(_03950_),
    .X(_04351_));
 sky130_fd_sc_hd__o211a_1 _11635_ (.A1(_03900_),
    .A2(_04343_),
    .B1(_04351_),
    .C1(_03954_),
    .X(_04352_));
 sky130_fd_sc_hd__mux2_1 _11636_ (.A0(\rbzero.tex_g0[43] ),
    .A1(\rbzero.tex_g0[42] ),
    .S(_04000_),
    .X(_04353_));
 sky130_fd_sc_hd__mux2_1 _11637_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_04000_),
    .X(_04354_));
 sky130_fd_sc_hd__mux2_1 _11638_ (.A0(_04353_),
    .A1(_04354_),
    .S(_04014_),
    .X(_04355_));
 sky130_fd_sc_hd__mux2_1 _11639_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(_04000_),
    .X(_04356_));
 sky130_fd_sc_hd__and2_1 _11640_ (.A(\rbzero.tex_g0[46] ),
    .B(_03925_),
    .X(_04357_));
 sky130_fd_sc_hd__a31o_1 _11641_ (.A1(\rbzero.tex_g0[47] ),
    .A2(_04142_),
    .A3(_04144_),
    .B1(_03915_),
    .X(_04358_));
 sky130_fd_sc_hd__o221a_1 _11642_ (.A1(_03957_),
    .A2(_04356_),
    .B1(_04357_),
    .B2(_04358_),
    .C1(_03920_),
    .X(_04359_));
 sky130_fd_sc_hd__a211o_1 _11643_ (.A1(_03972_),
    .A2(_04355_),
    .B1(_04359_),
    .C1(_03950_),
    .X(_04360_));
 sky130_fd_sc_hd__mux2_1 _11644_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_04000_),
    .X(_04361_));
 sky130_fd_sc_hd__mux2_1 _11645_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_04000_),
    .X(_04362_));
 sky130_fd_sc_hd__mux2_1 _11646_ (.A0(_04361_),
    .A1(_04362_),
    .S(_04014_),
    .X(_04363_));
 sky130_fd_sc_hd__mux2_1 _11647_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_04000_),
    .X(_04364_));
 sky130_fd_sc_hd__and3_1 _11648_ (.A(\rbzero.tex_g0[35] ),
    .B(_04142_),
    .C(_04144_),
    .X(_04365_));
 sky130_fd_sc_hd__a21o_1 _11649_ (.A1(\rbzero.tex_g0[34] ),
    .A2(_03961_),
    .B1(_03929_),
    .X(_04366_));
 sky130_fd_sc_hd__o221a_1 _11650_ (.A1(_03910_),
    .A2(_04364_),
    .B1(_04365_),
    .B2(_04366_),
    .C1(_03945_),
    .X(_04367_));
 sky130_fd_sc_hd__a211o_1 _11651_ (.A1(_03921_),
    .A2(_04363_),
    .B1(_04367_),
    .C1(_03899_),
    .X(_04368_));
 sky130_fd_sc_hd__a31o_1 _11652_ (.A1(_03985_),
    .A2(_04360_),
    .A3(_04368_),
    .B1(_03896_),
    .X(_04369_));
 sky130_fd_sc_hd__o32a_1 _11653_ (.A1(_04026_),
    .A2(_04318_),
    .A3(_04336_),
    .B1(_04352_),
    .B2(_04369_),
    .X(_04370_));
 sky130_fd_sc_hd__mux2_1 _11654_ (.A0(\rbzero.color_sky[2] ),
    .A1(\rbzero.color_floor[2] ),
    .S(_04030_),
    .X(_04371_));
 sky130_fd_sc_hd__mux2_1 _11655_ (.A0(_04370_),
    .A1(_04371_),
    .S(_04099_),
    .X(_04372_));
 sky130_fd_sc_hd__o21ba_1 _11656_ (.A1(_03826_),
    .A2(_04372_),
    .B1_N(_04117_),
    .X(_04373_));
 sky130_fd_sc_hd__buf_4 _11657_ (.A(_04373_),
    .X(o_rgb[14]));
 sky130_fd_sc_hd__clkbuf_4 _11658_ (.A(_03974_),
    .X(_04374_));
 sky130_fd_sc_hd__mux2_1 _11659_ (.A0(\rbzero.tex_g1[27] ),
    .A1(\rbzero.tex_g1[26] ),
    .S(_04374_),
    .X(_04375_));
 sky130_fd_sc_hd__mux2_1 _11660_ (.A0(\rbzero.tex_g1[25] ),
    .A1(\rbzero.tex_g1[24] ),
    .S(_04374_),
    .X(_04376_));
 sky130_fd_sc_hd__mux2_1 _11661_ (.A0(_04375_),
    .A1(_04376_),
    .S(_03968_),
    .X(_04377_));
 sky130_fd_sc_hd__clkbuf_4 _11662_ (.A(_03980_),
    .X(_04378_));
 sky130_fd_sc_hd__mux2_1 _11663_ (.A0(\rbzero.tex_g1[29] ),
    .A1(\rbzero.tex_g1[28] ),
    .S(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__and2_1 _11664_ (.A(\rbzero.tex_g1[30] ),
    .B(_04374_),
    .X(_04380_));
 sky130_fd_sc_hd__a31o_1 _11665_ (.A1(\rbzero.tex_g1[31] ),
    .A2(_03964_),
    .A3(_03965_),
    .B1(_03997_),
    .X(_04381_));
 sky130_fd_sc_hd__o221a_1 _11666_ (.A1(_03958_),
    .A2(_04379_),
    .B1(_04380_),
    .B2(_04381_),
    .C1(_04007_),
    .X(_04382_));
 sky130_fd_sc_hd__a211o_1 _11667_ (.A1(_03994_),
    .A2(_04377_),
    .B1(_04382_),
    .C1(_03956_),
    .X(_04383_));
 sky130_fd_sc_hd__mux2_1 _11668_ (.A0(\rbzero.tex_g1[19] ),
    .A1(\rbzero.tex_g1[18] ),
    .S(_04378_),
    .X(_04384_));
 sky130_fd_sc_hd__mux2_1 _11669_ (.A0(\rbzero.tex_g1[17] ),
    .A1(\rbzero.tex_g1[16] ),
    .S(_04378_),
    .X(_04385_));
 sky130_fd_sc_hd__mux2_1 _11670_ (.A0(_04384_),
    .A1(_04385_),
    .S(_03968_),
    .X(_04386_));
 sky130_fd_sc_hd__mux2_1 _11671_ (.A0(\rbzero.tex_g1[21] ),
    .A1(\rbzero.tex_g1[20] ),
    .S(_04378_),
    .X(_04387_));
 sky130_fd_sc_hd__and2_1 _11672_ (.A(\rbzero.tex_g1[22] ),
    .B(_04374_),
    .X(_04388_));
 sky130_fd_sc_hd__a31o_1 _11673_ (.A1(\rbzero.tex_g1[23] ),
    .A2(_03964_),
    .A3(_03965_),
    .B1(_03997_),
    .X(_04389_));
 sky130_fd_sc_hd__o221a_1 _11674_ (.A1(_03958_),
    .A2(_04387_),
    .B1(_04388_),
    .B2(_04389_),
    .C1(_04007_),
    .X(_04390_));
 sky130_fd_sc_hd__a211o_1 _11675_ (.A1(_03994_),
    .A2(_04386_),
    .B1(_04390_),
    .C1(_03900_),
    .X(_04391_));
 sky130_fd_sc_hd__and3_1 _11676_ (.A(\rbzero.tex_g1[3] ),
    .B(_03964_),
    .C(_03965_),
    .X(_04392_));
 sky130_fd_sc_hd__a21o_1 _11677_ (.A1(\rbzero.tex_g1[2] ),
    .A2(_04374_),
    .B1(_03997_),
    .X(_04393_));
 sky130_fd_sc_hd__mux2_1 _11678_ (.A0(\rbzero.tex_g1[1] ),
    .A1(\rbzero.tex_g1[0] ),
    .S(_03962_),
    .X(_04394_));
 sky130_fd_sc_hd__o221a_1 _11679_ (.A1(_04392_),
    .A2(_04393_),
    .B1(_04394_),
    .B2(_03958_),
    .C1(_03994_),
    .X(_04395_));
 sky130_fd_sc_hd__mux2_1 _11680_ (.A0(\rbzero.tex_g1[5] ),
    .A1(\rbzero.tex_g1[4] ),
    .S(_03962_),
    .X(_04396_));
 sky130_fd_sc_hd__and2_1 _11681_ (.A(\rbzero.tex_g1[6] ),
    .B(_04374_),
    .X(_04397_));
 sky130_fd_sc_hd__a31o_1 _11682_ (.A1(\rbzero.tex_g1[7] ),
    .A2(_03964_),
    .A3(_03965_),
    .B1(_03997_),
    .X(_04398_));
 sky130_fd_sc_hd__o221a_1 _11683_ (.A1(_03958_),
    .A2(_04396_),
    .B1(_04397_),
    .B2(_04398_),
    .C1(_04007_),
    .X(_04399_));
 sky130_fd_sc_hd__mux2_1 _11684_ (.A0(\rbzero.tex_g1[15] ),
    .A1(\rbzero.tex_g1[14] ),
    .S(_03980_),
    .X(_04400_));
 sky130_fd_sc_hd__mux2_1 _11685_ (.A0(\rbzero.tex_g1[13] ),
    .A1(\rbzero.tex_g1[12] ),
    .S(_03980_),
    .X(_04401_));
 sky130_fd_sc_hd__mux2_1 _11686_ (.A0(_04400_),
    .A1(_04401_),
    .S(_03997_),
    .X(_04402_));
 sky130_fd_sc_hd__mux2_1 _11687_ (.A0(\rbzero.tex_g1[9] ),
    .A1(\rbzero.tex_g1[8] ),
    .S(_03980_),
    .X(_04403_));
 sky130_fd_sc_hd__and3_1 _11688_ (.A(\rbzero.tex_g1[11] ),
    .B(_04143_),
    .C(_04145_),
    .X(_04404_));
 sky130_fd_sc_hd__a21o_1 _11689_ (.A1(\rbzero.tex_g1[10] ),
    .A2(_03959_),
    .B1(_03916_),
    .X(_04405_));
 sky130_fd_sc_hd__o221a_1 _11690_ (.A1(_04323_),
    .A2(_04403_),
    .B1(_04404_),
    .B2(_04405_),
    .C1(_03972_),
    .X(_04406_));
 sky130_fd_sc_hd__a211o_1 _11691_ (.A1(_04007_),
    .A2(_04402_),
    .B1(_04406_),
    .C1(_03956_),
    .X(_04407_));
 sky130_fd_sc_hd__o311a_1 _11692_ (.A1(_03900_),
    .A2(_04395_),
    .A3(_04399_),
    .B1(_03985_),
    .C1(_04407_),
    .X(_04408_));
 sky130_fd_sc_hd__a311o_1 _11693_ (.A1(_03954_),
    .A2(_04383_),
    .A3(_04391_),
    .B1(_04408_),
    .C1(_04026_),
    .X(_04409_));
 sky130_fd_sc_hd__mux2_1 _11694_ (.A0(\rbzero.tex_g1[63] ),
    .A1(\rbzero.tex_g1[62] ),
    .S(_04378_),
    .X(_04410_));
 sky130_fd_sc_hd__mux2_1 _11695_ (.A0(\rbzero.tex_g1[61] ),
    .A1(\rbzero.tex_g1[60] ),
    .S(_04378_),
    .X(_04411_));
 sky130_fd_sc_hd__mux2_1 _11696_ (.A0(_04410_),
    .A1(_04411_),
    .S(_03968_),
    .X(_04412_));
 sky130_fd_sc_hd__mux2_1 _11697_ (.A0(\rbzero.tex_g1[57] ),
    .A1(\rbzero.tex_g1[56] ),
    .S(_04378_),
    .X(_04413_));
 sky130_fd_sc_hd__and2_1 _11698_ (.A(\rbzero.tex_g1[58] ),
    .B(_04374_),
    .X(_04414_));
 sky130_fd_sc_hd__a31o_1 _11699_ (.A1(\rbzero.tex_g1[59] ),
    .A2(_03964_),
    .A3(_03965_),
    .B1(_03997_),
    .X(_04415_));
 sky130_fd_sc_hd__o221a_1 _11700_ (.A1(_03958_),
    .A2(_04413_),
    .B1(_04414_),
    .B2(_04415_),
    .C1(_03994_),
    .X(_04416_));
 sky130_fd_sc_hd__a211o_1 _11701_ (.A1(_04007_),
    .A2(_04412_),
    .B1(_04416_),
    .C1(_03956_),
    .X(_04417_));
 sky130_fd_sc_hd__mux2_1 _11702_ (.A0(\rbzero.tex_g1[49] ),
    .A1(\rbzero.tex_g1[48] ),
    .S(_04378_),
    .X(_04418_));
 sky130_fd_sc_hd__mux2_1 _11703_ (.A0(\rbzero.tex_g1[51] ),
    .A1(\rbzero.tex_g1[50] ),
    .S(_04378_),
    .X(_04419_));
 sky130_fd_sc_hd__mux2_1 _11704_ (.A0(_04418_),
    .A1(_04419_),
    .S(_03958_),
    .X(_04420_));
 sky130_fd_sc_hd__and2_1 _11705_ (.A(\rbzero.tex_g1[54] ),
    .B(_04374_),
    .X(_04421_));
 sky130_fd_sc_hd__a31o_1 _11706_ (.A1(\rbzero.tex_g1[55] ),
    .A2(_03964_),
    .A3(_03965_),
    .B1(_03997_),
    .X(_04422_));
 sky130_fd_sc_hd__mux2_1 _11707_ (.A0(\rbzero.tex_g1[53] ),
    .A1(\rbzero.tex_g1[52] ),
    .S(_04378_),
    .X(_04423_));
 sky130_fd_sc_hd__o221a_1 _11708_ (.A1(_04421_),
    .A2(_04422_),
    .B1(_04423_),
    .B2(_03958_),
    .C1(_04007_),
    .X(_04424_));
 sky130_fd_sc_hd__a211o_1 _11709_ (.A1(_03994_),
    .A2(_04420_),
    .B1(_04424_),
    .C1(_03900_),
    .X(_04425_));
 sky130_fd_sc_hd__mux2_1 _11710_ (.A0(\rbzero.tex_g1[45] ),
    .A1(\rbzero.tex_g1[44] ),
    .S(_03962_),
    .X(_04426_));
 sky130_fd_sc_hd__and2_1 _11711_ (.A(\rbzero.tex_g1[46] ),
    .B(_04374_),
    .X(_04427_));
 sky130_fd_sc_hd__a31o_1 _11712_ (.A1(\rbzero.tex_g1[47] ),
    .A2(_03964_),
    .A3(_03965_),
    .B1(_03997_),
    .X(_04428_));
 sky130_fd_sc_hd__o221a_1 _11713_ (.A1(_03958_),
    .A2(_04426_),
    .B1(_04427_),
    .B2(_04428_),
    .C1(_03924_),
    .X(_04429_));
 sky130_fd_sc_hd__mux2_1 _11714_ (.A0(\rbzero.tex_g1[43] ),
    .A1(\rbzero.tex_g1[42] ),
    .S(_03962_),
    .X(_04430_));
 sky130_fd_sc_hd__and2_1 _11715_ (.A(\rbzero.tex_g1[40] ),
    .B(_04374_),
    .X(_04431_));
 sky130_fd_sc_hd__a31o_1 _11716_ (.A1(\rbzero.tex_g1[41] ),
    .A2(_03964_),
    .A3(_03965_),
    .B1(_03932_),
    .X(_04432_));
 sky130_fd_sc_hd__o221a_1 _11717_ (.A1(_03968_),
    .A2(_04430_),
    .B1(_04431_),
    .B2(_04432_),
    .C1(_03994_),
    .X(_04433_));
 sky130_fd_sc_hd__mux2_1 _11718_ (.A0(\rbzero.tex_g1[39] ),
    .A1(\rbzero.tex_g1[38] ),
    .S(_03980_),
    .X(_04434_));
 sky130_fd_sc_hd__mux2_1 _11719_ (.A0(\rbzero.tex_g1[37] ),
    .A1(\rbzero.tex_g1[36] ),
    .S(_03980_),
    .X(_04435_));
 sky130_fd_sc_hd__mux2_1 _11720_ (.A0(_04434_),
    .A1(_04435_),
    .S(_03997_),
    .X(_04436_));
 sky130_fd_sc_hd__mux2_1 _11721_ (.A0(\rbzero.tex_g1[33] ),
    .A1(\rbzero.tex_g1[32] ),
    .S(_03980_),
    .X(_04437_));
 sky130_fd_sc_hd__and3_1 _11722_ (.A(\rbzero.tex_g1[35] ),
    .B(_03939_),
    .C(_03941_),
    .X(_04438_));
 sky130_fd_sc_hd__a21o_1 _11723_ (.A1(\rbzero.tex_g1[34] ),
    .A2(_03959_),
    .B1(_03916_),
    .X(_04439_));
 sky130_fd_sc_hd__o221a_1 _11724_ (.A1(_04323_),
    .A2(_04437_),
    .B1(_04438_),
    .B2(_04439_),
    .C1(_03972_),
    .X(_04440_));
 sky130_fd_sc_hd__a211o_1 _11725_ (.A1(_04007_),
    .A2(_04436_),
    .B1(_04440_),
    .C1(_03899_),
    .X(_04441_));
 sky130_fd_sc_hd__o311a_1 _11726_ (.A1(_03956_),
    .A2(_04429_),
    .A3(_04433_),
    .B1(_04441_),
    .C1(_03985_),
    .X(_04442_));
 sky130_fd_sc_hd__a311o_1 _11727_ (.A1(_03954_),
    .A2(_04417_),
    .A3(_04425_),
    .B1(_04442_),
    .C1(_03896_),
    .X(_04443_));
 sky130_fd_sc_hd__nand3b_2 _11728_ (.A_N(_04099_),
    .B(_04409_),
    .C(_04443_),
    .Y(_04444_));
 sky130_fd_sc_hd__mux2_1 _11729_ (.A0(\rbzero.color_sky[3] ),
    .A1(\rbzero.color_floor[3] ),
    .S(_04030_),
    .X(_04445_));
 sky130_fd_sc_hd__nand2_1 _11730_ (.A(_04099_),
    .B(_04445_),
    .Y(_04446_));
 sky130_fd_sc_hd__a31o_4 _11731_ (.A1(_03825_),
    .A2(_04444_),
    .A3(_04446_),
    .B1(_04301_),
    .X(_04447_));
 sky130_fd_sc_hd__inv_2 _11732_ (.A(_04447_),
    .Y(o_rgb[15]));
 sky130_fd_sc_hd__mux2_1 _11733_ (.A0(\rbzero.tex_b0[63] ),
    .A1(\rbzero.tex_b0[62] ),
    .S(_04013_),
    .X(_04448_));
 sky130_fd_sc_hd__mux2_1 _11734_ (.A0(\rbzero.tex_b0[61] ),
    .A1(\rbzero.tex_b0[60] ),
    .S(_04013_),
    .X(_04449_));
 sky130_fd_sc_hd__mux2_1 _11735_ (.A0(_04448_),
    .A1(_04449_),
    .S(_03968_),
    .X(_04450_));
 sky130_fd_sc_hd__mux2_1 _11736_ (.A0(\rbzero.tex_b0[57] ),
    .A1(\rbzero.tex_b0[56] ),
    .S(_04013_),
    .X(_04451_));
 sky130_fd_sc_hd__and2_1 _11737_ (.A(\rbzero.tex_b0[58] ),
    .B(_03962_),
    .X(_04452_));
 sky130_fd_sc_hd__a31o_1 _11738_ (.A1(\rbzero.tex_b0[59] ),
    .A2(_04143_),
    .A3(_04145_),
    .B1(_03930_),
    .X(_04453_));
 sky130_fd_sc_hd__o221a_1 _11739_ (.A1(_04323_),
    .A2(_04451_),
    .B1(_04452_),
    .B2(_04453_),
    .C1(_03972_),
    .X(_04454_));
 sky130_fd_sc_hd__a211o_1 _11740_ (.A1(_04007_),
    .A2(_04450_),
    .B1(_04454_),
    .C1(_03956_),
    .X(_04455_));
 sky130_fd_sc_hd__mux2_1 _11741_ (.A0(\rbzero.tex_b0[49] ),
    .A1(\rbzero.tex_b0[48] ),
    .S(_04013_),
    .X(_04456_));
 sky130_fd_sc_hd__mux2_1 _11742_ (.A0(\rbzero.tex_b0[51] ),
    .A1(\rbzero.tex_b0[50] ),
    .S(_04013_),
    .X(_04457_));
 sky130_fd_sc_hd__mux2_1 _11743_ (.A0(_04456_),
    .A1(_04457_),
    .S(_04323_),
    .X(_04458_));
 sky130_fd_sc_hd__and2_1 _11744_ (.A(\rbzero.tex_b0[54] ),
    .B(_03959_),
    .X(_04459_));
 sky130_fd_sc_hd__a31o_1 _11745_ (.A1(\rbzero.tex_b0[55] ),
    .A2(_04143_),
    .A3(_04145_),
    .B1(_03930_),
    .X(_04460_));
 sky130_fd_sc_hd__mux2_1 _11746_ (.A0(\rbzero.tex_b0[53] ),
    .A1(\rbzero.tex_b0[52] ),
    .S(_03959_),
    .X(_04461_));
 sky130_fd_sc_hd__o221a_1 _11747_ (.A1(_04459_),
    .A2(_04460_),
    .B1(_04461_),
    .B2(_03958_),
    .C1(_03924_),
    .X(_04462_));
 sky130_fd_sc_hd__a211o_1 _11748_ (.A1(_03994_),
    .A2(_04458_),
    .B1(_04462_),
    .C1(_03900_),
    .X(_04463_));
 sky130_fd_sc_hd__mux2_1 _11749_ (.A0(\rbzero.tex_b0[45] ),
    .A1(\rbzero.tex_b0[44] ),
    .S(_03980_),
    .X(_04464_));
 sky130_fd_sc_hd__and2_1 _11750_ (.A(\rbzero.tex_b0[46] ),
    .B(_03959_),
    .X(_04465_));
 sky130_fd_sc_hd__a31o_1 _11751_ (.A1(\rbzero.tex_b0[47] ),
    .A2(_04143_),
    .A3(_04145_),
    .B1(_03916_),
    .X(_04466_));
 sky130_fd_sc_hd__o221a_1 _11752_ (.A1(_04323_),
    .A2(_04464_),
    .B1(_04465_),
    .B2(_04466_),
    .C1(_03921_),
    .X(_04467_));
 sky130_fd_sc_hd__mux2_1 _11753_ (.A0(\rbzero.tex_b0[43] ),
    .A1(\rbzero.tex_b0[42] ),
    .S(_04001_),
    .X(_04468_));
 sky130_fd_sc_hd__and2_1 _11754_ (.A(\rbzero.tex_b0[40] ),
    .B(_03962_),
    .X(_04469_));
 sky130_fd_sc_hd__a31o_1 _11755_ (.A1(\rbzero.tex_b0[41] ),
    .A2(_04143_),
    .A3(_04145_),
    .B1(_03957_),
    .X(_04470_));
 sky130_fd_sc_hd__o221a_1 _11756_ (.A1(_03968_),
    .A2(_04468_),
    .B1(_04469_),
    .B2(_04470_),
    .C1(_03972_),
    .X(_04471_));
 sky130_fd_sc_hd__mux2_1 _11757_ (.A0(\rbzero.tex_b0[39] ),
    .A1(\rbzero.tex_b0[38] ),
    .S(_03904_),
    .X(_04472_));
 sky130_fd_sc_hd__mux2_1 _11758_ (.A0(\rbzero.tex_b0[37] ),
    .A1(\rbzero.tex_b0[36] ),
    .S(_03904_),
    .X(_04473_));
 sky130_fd_sc_hd__mux2_1 _11759_ (.A0(_04472_),
    .A1(_04473_),
    .S(_03916_),
    .X(_04474_));
 sky130_fd_sc_hd__mux2_1 _11760_ (.A0(\rbzero.tex_b0[33] ),
    .A1(\rbzero.tex_b0[32] ),
    .S(_03904_),
    .X(_04475_));
 sky130_fd_sc_hd__and3_1 _11761_ (.A(\rbzero.tex_b0[35] ),
    .B(_04142_),
    .C(_04144_),
    .X(_04476_));
 sky130_fd_sc_hd__a21o_1 _11762_ (.A1(\rbzero.tex_b0[34] ),
    .A2(_03936_),
    .B1(_03929_),
    .X(_04477_));
 sky130_fd_sc_hd__o221a_1 _11763_ (.A1(_03957_),
    .A2(_04475_),
    .B1(_04476_),
    .B2(_04477_),
    .C1(_03946_),
    .X(_04478_));
 sky130_fd_sc_hd__a211o_1 _11764_ (.A1(_03924_),
    .A2(_04474_),
    .B1(_04478_),
    .C1(_03899_),
    .X(_04479_));
 sky130_fd_sc_hd__o311a_1 _11765_ (.A1(_03956_),
    .A2(_04467_),
    .A3(_04471_),
    .B1(_04479_),
    .C1(_03985_),
    .X(_04480_));
 sky130_fd_sc_hd__a311o_1 _11766_ (.A1(_03954_),
    .A2(_04455_),
    .A3(_04463_),
    .B1(_04480_),
    .C1(_03896_),
    .X(_04481_));
 sky130_fd_sc_hd__mux2_1 _11767_ (.A0(\rbzero.tex_b0[27] ),
    .A1(\rbzero.tex_b0[26] ),
    .S(_04013_),
    .X(_04482_));
 sky130_fd_sc_hd__mux2_1 _11768_ (.A0(\rbzero.tex_b0[25] ),
    .A1(\rbzero.tex_b0[24] ),
    .S(_04001_),
    .X(_04483_));
 sky130_fd_sc_hd__mux2_1 _11769_ (.A0(_04482_),
    .A1(_04483_),
    .S(_03968_),
    .X(_04484_));
 sky130_fd_sc_hd__mux2_1 _11770_ (.A0(\rbzero.tex_b0[29] ),
    .A1(\rbzero.tex_b0[28] ),
    .S(_04001_),
    .X(_04485_));
 sky130_fd_sc_hd__and2_1 _11771_ (.A(\rbzero.tex_b0[30] ),
    .B(_03962_),
    .X(_04486_));
 sky130_fd_sc_hd__a31o_1 _11772_ (.A1(\rbzero.tex_b0[31] ),
    .A2(_04143_),
    .A3(_04145_),
    .B1(_03930_),
    .X(_04487_));
 sky130_fd_sc_hd__o221a_1 _11773_ (.A1(_04323_),
    .A2(_04485_),
    .B1(_04486_),
    .B2(_04487_),
    .C1(_03921_),
    .X(_04488_));
 sky130_fd_sc_hd__a211o_1 _11774_ (.A1(_03994_),
    .A2(_04484_),
    .B1(_04488_),
    .C1(_03956_),
    .X(_04489_));
 sky130_fd_sc_hd__mux2_1 _11775_ (.A0(\rbzero.tex_b0[19] ),
    .A1(\rbzero.tex_b0[18] ),
    .S(_04001_),
    .X(_04490_));
 sky130_fd_sc_hd__mux2_1 _11776_ (.A0(\rbzero.tex_b0[17] ),
    .A1(\rbzero.tex_b0[16] ),
    .S(_04001_),
    .X(_04491_));
 sky130_fd_sc_hd__mux2_1 _11777_ (.A0(_04490_),
    .A1(_04491_),
    .S(_03968_),
    .X(_04492_));
 sky130_fd_sc_hd__mux2_1 _11778_ (.A0(\rbzero.tex_b0[21] ),
    .A1(\rbzero.tex_b0[20] ),
    .S(_04001_),
    .X(_04493_));
 sky130_fd_sc_hd__and2_1 _11779_ (.A(\rbzero.tex_b0[22] ),
    .B(_03962_),
    .X(_04494_));
 sky130_fd_sc_hd__a31o_1 _11780_ (.A1(\rbzero.tex_b0[23] ),
    .A2(_04143_),
    .A3(_04145_),
    .B1(_03930_),
    .X(_04495_));
 sky130_fd_sc_hd__o221a_1 _11781_ (.A1(_04323_),
    .A2(_04493_),
    .B1(_04494_),
    .B2(_04495_),
    .C1(_03921_),
    .X(_04496_));
 sky130_fd_sc_hd__a211o_1 _11782_ (.A1(_03994_),
    .A2(_04492_),
    .B1(_04496_),
    .C1(_03900_),
    .X(_04497_));
 sky130_fd_sc_hd__and3_1 _11783_ (.A(\rbzero.tex_b0[3] ),
    .B(_04143_),
    .C(_04145_),
    .X(_04498_));
 sky130_fd_sc_hd__a21o_1 _11784_ (.A1(\rbzero.tex_b0[2] ),
    .A2(_03959_),
    .B1(_03916_),
    .X(_04499_));
 sky130_fd_sc_hd__mux2_1 _11785_ (.A0(\rbzero.tex_b0[1] ),
    .A1(\rbzero.tex_b0[0] ),
    .S(_04001_),
    .X(_04500_));
 sky130_fd_sc_hd__o221a_1 _11786_ (.A1(_04498_),
    .A2(_04499_),
    .B1(_04500_),
    .B2(_04323_),
    .C1(_03972_),
    .X(_04501_));
 sky130_fd_sc_hd__mux2_1 _11787_ (.A0(\rbzero.tex_b0[5] ),
    .A1(\rbzero.tex_b0[4] ),
    .S(_04001_),
    .X(_04502_));
 sky130_fd_sc_hd__and2_1 _11788_ (.A(\rbzero.tex_b0[6] ),
    .B(_03959_),
    .X(_04503_));
 sky130_fd_sc_hd__a31o_1 _11789_ (.A1(\rbzero.tex_b0[7] ),
    .A2(_04143_),
    .A3(_04145_),
    .B1(_03930_),
    .X(_04504_));
 sky130_fd_sc_hd__o221a_1 _11790_ (.A1(_04323_),
    .A2(_04502_),
    .B1(_04503_),
    .B2(_04504_),
    .C1(_03921_),
    .X(_04505_));
 sky130_fd_sc_hd__mux2_1 _11791_ (.A0(\rbzero.tex_b0[15] ),
    .A1(\rbzero.tex_b0[14] ),
    .S(_03925_),
    .X(_04506_));
 sky130_fd_sc_hd__mux2_1 _11792_ (.A0(\rbzero.tex_b0[13] ),
    .A1(\rbzero.tex_b0[12] ),
    .S(_03925_),
    .X(_04507_));
 sky130_fd_sc_hd__mux2_1 _11793_ (.A0(_04506_),
    .A1(_04507_),
    .S(_03916_),
    .X(_04508_));
 sky130_fd_sc_hd__mux2_1 _11794_ (.A0(\rbzero.tex_b0[9] ),
    .A1(\rbzero.tex_b0[8] ),
    .S(_03925_),
    .X(_04509_));
 sky130_fd_sc_hd__and3_1 _11795_ (.A(\rbzero.tex_b0[11] ),
    .B(_04142_),
    .C(_04144_),
    .X(_04510_));
 sky130_fd_sc_hd__a21o_1 _11796_ (.A1(\rbzero.tex_b0[10] ),
    .A2(_03936_),
    .B1(_03929_),
    .X(_04511_));
 sky130_fd_sc_hd__o221a_1 _11797_ (.A1(_03957_),
    .A2(_04509_),
    .B1(_04510_),
    .B2(_04511_),
    .C1(_03946_),
    .X(_04512_));
 sky130_fd_sc_hd__a211o_1 _11798_ (.A1(_03924_),
    .A2(_04508_),
    .B1(_04512_),
    .C1(_03950_),
    .X(_04513_));
 sky130_fd_sc_hd__o311a_1 _11799_ (.A1(_03900_),
    .A2(_04501_),
    .A3(_04505_),
    .B1(_03985_),
    .C1(_04513_),
    .X(_04514_));
 sky130_fd_sc_hd__a311o_1 _11800_ (.A1(_03954_),
    .A2(_04489_),
    .A3(_04497_),
    .B1(_04514_),
    .C1(_04026_),
    .X(_04515_));
 sky130_fd_sc_hd__nand3b_2 _11801_ (.A_N(_04099_),
    .B(_04481_),
    .C(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hd__mux2_1 _11802_ (.A0(\rbzero.color_sky[4] ),
    .A1(\rbzero.color_floor[4] ),
    .S(_04030_),
    .X(_04517_));
 sky130_fd_sc_hd__nand2_1 _11803_ (.A(_04099_),
    .B(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__a31o_4 _11804_ (.A1(_03825_),
    .A2(_04516_),
    .A3(_04518_),
    .B1(_04117_),
    .X(_04519_));
 sky130_fd_sc_hd__inv_2 _11805_ (.A(_04519_),
    .Y(o_rgb[22]));
 sky130_fd_sc_hd__mux2_1 _11806_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(_04032_),
    .X(_04520_));
 sky130_fd_sc_hd__mux2_1 _11807_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_04032_),
    .X(_04521_));
 sky130_fd_sc_hd__mux2_1 _11808_ (.A0(_04520_),
    .A1(_04521_),
    .S(_03908_),
    .X(_04522_));
 sky130_fd_sc_hd__mux2_1 _11809_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(_04032_),
    .X(_04523_));
 sky130_fd_sc_hd__mux2_1 _11810_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(_04032_),
    .X(_04524_));
 sky130_fd_sc_hd__mux2_1 _11811_ (.A0(_04523_),
    .A1(_04524_),
    .S(_03928_),
    .X(_04525_));
 sky130_fd_sc_hd__mux2_1 _11812_ (.A0(_04522_),
    .A1(_04525_),
    .S(_03919_),
    .X(_04526_));
 sky130_fd_sc_hd__mux2_1 _11813_ (.A0(\rbzero.tex_b1[63] ),
    .A1(\rbzero.tex_b1[62] ),
    .S(_04032_),
    .X(_04527_));
 sky130_fd_sc_hd__mux2_1 _11814_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_04032_),
    .X(_04528_));
 sky130_fd_sc_hd__mux2_1 _11815_ (.A0(_04527_),
    .A1(_04528_),
    .S(_03928_),
    .X(_04529_));
 sky130_fd_sc_hd__mux2_1 _11816_ (.A0(\rbzero.tex_b1[57] ),
    .A1(\rbzero.tex_b1[56] ),
    .S(_04032_),
    .X(_04530_));
 sky130_fd_sc_hd__and2_1 _11817_ (.A(\rbzero.tex_b1[58] ),
    .B(_03934_),
    .X(_04531_));
 sky130_fd_sc_hd__a31o_1 _11818_ (.A1(\rbzero.tex_b1[59] ),
    .A2(_03859_),
    .A3(_03901_),
    .B1(_03914_),
    .X(_04532_));
 sky130_fd_sc_hd__o221a_1 _11819_ (.A1(_03908_),
    .A2(_04530_),
    .B1(_04531_),
    .B2(_04532_),
    .C1(_03944_),
    .X(_04533_));
 sky130_fd_sc_hd__a211o_1 _11820_ (.A1(_03920_),
    .A2(_04529_),
    .B1(_04533_),
    .C1(_03949_),
    .X(_04534_));
 sky130_fd_sc_hd__o211a_1 _11821_ (.A1(_03898_),
    .A2(_04526_),
    .B1(_04534_),
    .C1(_03953_),
    .X(_04535_));
 sky130_fd_sc_hd__mux2_1 _11822_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(_03903_),
    .X(_04536_));
 sky130_fd_sc_hd__and2_1 _11823_ (.A(\rbzero.tex_b1[46] ),
    .B(_04119_),
    .X(_04537_));
 sky130_fd_sc_hd__a31o_1 _11824_ (.A1(\rbzero.tex_b1[47] ),
    .A2(_03938_),
    .A3(_03940_),
    .B1(_03915_),
    .X(_04538_));
 sky130_fd_sc_hd__o221a_1 _11825_ (.A1(_03909_),
    .A2(_04536_),
    .B1(_04537_),
    .B2(_04538_),
    .C1(_03920_),
    .X(_04539_));
 sky130_fd_sc_hd__mux2_1 _11826_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(_03903_),
    .X(_04540_));
 sky130_fd_sc_hd__and2_1 _11827_ (.A(\rbzero.tex_b1[40] ),
    .B(_04119_),
    .X(_04541_));
 sky130_fd_sc_hd__a31o_1 _11828_ (.A1(\rbzero.tex_b1[41] ),
    .A2(_03938_),
    .A3(_03940_),
    .B1(_03908_),
    .X(_04542_));
 sky130_fd_sc_hd__o221a_1 _11829_ (.A1(_03929_),
    .A2(_04540_),
    .B1(_04541_),
    .B2(_04542_),
    .C1(_03945_),
    .X(_04543_));
 sky130_fd_sc_hd__clkbuf_4 _11830_ (.A(_03902_),
    .X(_04544_));
 sky130_fd_sc_hd__mux2_1 _11831_ (.A0(\rbzero.tex_b1[39] ),
    .A1(\rbzero.tex_b1[38] ),
    .S(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__mux2_1 _11832_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(_04032_),
    .X(_04546_));
 sky130_fd_sc_hd__mux2_1 _11833_ (.A0(_04545_),
    .A1(_04546_),
    .S(_03928_),
    .X(_04547_));
 sky130_fd_sc_hd__mux2_1 _11834_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(_04032_),
    .X(_04548_));
 sky130_fd_sc_hd__and3_1 _11835_ (.A(\rbzero.tex_b1[35] ),
    .B(_03859_),
    .C(_03901_),
    .X(_04549_));
 sky130_fd_sc_hd__a21o_1 _11836_ (.A1(\rbzero.tex_b1[34] ),
    .A2(_03934_),
    .B1(_03928_),
    .X(_04550_));
 sky130_fd_sc_hd__o221a_1 _11837_ (.A1(_03908_),
    .A2(_04548_),
    .B1(_04549_),
    .B2(_04550_),
    .C1(_03944_),
    .X(_04551_));
 sky130_fd_sc_hd__a211o_1 _11838_ (.A1(_03920_),
    .A2(_04547_),
    .B1(_04551_),
    .C1(_03898_),
    .X(_04552_));
 sky130_fd_sc_hd__o311a_1 _11839_ (.A1(_03949_),
    .A2(_04539_),
    .A3(_04543_),
    .B1(_04552_),
    .C1(_03984_),
    .X(_04553_));
 sky130_fd_sc_hd__mux2_1 _11840_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(_04544_),
    .X(_04554_));
 sky130_fd_sc_hd__mux2_1 _11841_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(_04544_),
    .X(_04555_));
 sky130_fd_sc_hd__mux2_1 _11842_ (.A0(_04554_),
    .A1(_04555_),
    .S(_03928_),
    .X(_04556_));
 sky130_fd_sc_hd__mux2_1 _11843_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(_04544_),
    .X(_04557_));
 sky130_fd_sc_hd__mux2_1 _11844_ (.A0(\rbzero.tex_b1[23] ),
    .A1(\rbzero.tex_b1[22] ),
    .S(_04544_),
    .X(_04558_));
 sky130_fd_sc_hd__mux2_1 _11845_ (.A0(_04557_),
    .A1(_04558_),
    .S(_03908_),
    .X(_04559_));
 sky130_fd_sc_hd__mux2_1 _11846_ (.A0(_04556_),
    .A1(_04559_),
    .S(_03920_),
    .X(_04560_));
 sky130_fd_sc_hd__mux2_1 _11847_ (.A0(\rbzero.tex_b1[27] ),
    .A1(\rbzero.tex_b1[26] ),
    .S(_03934_),
    .X(_04561_));
 sky130_fd_sc_hd__mux2_1 _11848_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(_03934_),
    .X(_04562_));
 sky130_fd_sc_hd__mux2_1 _11849_ (.A0(_04561_),
    .A1(_04562_),
    .S(_03915_),
    .X(_04563_));
 sky130_fd_sc_hd__mux2_1 _11850_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(_03934_),
    .X(_04564_));
 sky130_fd_sc_hd__and2_1 _11851_ (.A(\rbzero.tex_b1[30] ),
    .B(_03934_),
    .X(_04565_));
 sky130_fd_sc_hd__a31o_1 _11852_ (.A1(\rbzero.tex_b1[31] ),
    .A2(_03938_),
    .A3(_03940_),
    .B1(_03928_),
    .X(_04566_));
 sky130_fd_sc_hd__o221a_1 _11853_ (.A1(_03909_),
    .A2(_04564_),
    .B1(_04565_),
    .B2(_04566_),
    .C1(_03919_),
    .X(_04567_));
 sky130_fd_sc_hd__a211o_1 _11854_ (.A1(_03945_),
    .A2(_04563_),
    .B1(_04567_),
    .C1(_03949_),
    .X(_04568_));
 sky130_fd_sc_hd__o211a_1 _11855_ (.A1(_03898_),
    .A2(_04560_),
    .B1(_04568_),
    .C1(_03953_),
    .X(_04569_));
 sky130_fd_sc_hd__mux2_1 _11856_ (.A0(\rbzero.tex_b1[15] ),
    .A1(\rbzero.tex_b1[14] ),
    .S(_04544_),
    .X(_04570_));
 sky130_fd_sc_hd__mux2_1 _11857_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_04544_),
    .X(_04571_));
 sky130_fd_sc_hd__mux2_1 _11858_ (.A0(_04570_),
    .A1(_04571_),
    .S(_03915_),
    .X(_04572_));
 sky130_fd_sc_hd__mux2_1 _11859_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_04544_),
    .X(_04573_));
 sky130_fd_sc_hd__and3_1 _11860_ (.A(\rbzero.tex_b1[11] ),
    .B(_03938_),
    .C(_03940_),
    .X(_04574_));
 sky130_fd_sc_hd__a21o_1 _11861_ (.A1(\rbzero.tex_b1[10] ),
    .A2(_03903_),
    .B1(_03928_),
    .X(_04575_));
 sky130_fd_sc_hd__o221a_1 _11862_ (.A1(_03909_),
    .A2(_04573_),
    .B1(_04574_),
    .B2(_04575_),
    .C1(_03944_),
    .X(_04576_));
 sky130_fd_sc_hd__a211o_1 _11863_ (.A1(_03920_),
    .A2(_04572_),
    .B1(_04576_),
    .C1(_03949_),
    .X(_04577_));
 sky130_fd_sc_hd__mux2_1 _11864_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_04544_),
    .X(_04578_));
 sky130_fd_sc_hd__mux2_1 _11865_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(_04544_),
    .X(_04579_));
 sky130_fd_sc_hd__mux2_1 _11866_ (.A0(_04578_),
    .A1(_04579_),
    .S(_03908_),
    .X(_04580_));
 sky130_fd_sc_hd__and3_1 _11867_ (.A(\rbzero.tex_b1[3] ),
    .B(_03859_),
    .C(_03901_),
    .X(_04581_));
 sky130_fd_sc_hd__a21o_1 _11868_ (.A1(\rbzero.tex_b1[2] ),
    .A2(_03903_),
    .B1(_03928_),
    .X(_04582_));
 sky130_fd_sc_hd__mux2_1 _11869_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[0] ),
    .S(_03934_),
    .X(_04583_));
 sky130_fd_sc_hd__o221a_1 _11870_ (.A1(_04581_),
    .A2(_04582_),
    .B1(_04583_),
    .B2(_03909_),
    .C1(_03944_),
    .X(_04584_));
 sky130_fd_sc_hd__a211o_1 _11871_ (.A1(_03920_),
    .A2(_04580_),
    .B1(_04584_),
    .C1(_03898_),
    .X(_04585_));
 sky130_fd_sc_hd__a31o_1 _11872_ (.A1(_03984_),
    .A2(_04577_),
    .A3(_04585_),
    .B1(_04026_),
    .X(_04586_));
 sky130_fd_sc_hd__o32a_1 _11873_ (.A1(_03896_),
    .A2(_04535_),
    .A3(_04553_),
    .B1(_04569_),
    .B2(_04586_),
    .X(_04587_));
 sky130_fd_sc_hd__mux2_1 _11874_ (.A0(\rbzero.color_sky[5] ),
    .A1(\rbzero.color_floor[5] ),
    .S(_04030_),
    .X(_04588_));
 sky130_fd_sc_hd__mux2_1 _11875_ (.A0(_04587_),
    .A1(_04588_),
    .S(_04099_),
    .X(_04589_));
 sky130_fd_sc_hd__o21ba_1 _11876_ (.A1(_03826_),
    .A2(_04589_),
    .B1_N(_04301_),
    .X(_04590_));
 sky130_fd_sc_hd__buf_4 _11877_ (.A(_04590_),
    .X(o_rgb[23]));
 sky130_fd_sc_hd__buf_2 _11878_ (.A(\gpout0.hpos[2] ),
    .X(_04591_));
 sky130_fd_sc_hd__clkbuf_4 _11879_ (.A(\gpout0.hpos[1] ),
    .X(_04592_));
 sky130_fd_sc_hd__nand2_1 _11880_ (.A(_04592_),
    .B(_03289_),
    .Y(_04593_));
 sky130_fd_sc_hd__o21a_1 _11881_ (.A1(_04592_),
    .A2(\rbzero.row_render.wall[1] ),
    .B1(_03288_),
    .X(_04594_));
 sky130_fd_sc_hd__inv_2 _11882_ (.A(\rbzero.row_render.wall[0] ),
    .Y(_04595_));
 sky130_fd_sc_hd__inv_2 _11883_ (.A(\rbzero.row_render.wall[1] ),
    .Y(_04596_));
 sky130_fd_sc_hd__a211o_1 _11884_ (.A1(_03288_),
    .A2(_04596_),
    .B1(\rbzero.row_render.wall[0] ),
    .C1(_04592_),
    .X(_04597_));
 sky130_fd_sc_hd__o221a_1 _11885_ (.A1(\rbzero.row_render.side ),
    .A2(_04593_),
    .B1(_04594_),
    .B2(_04595_),
    .C1(_04597_),
    .X(_04598_));
 sky130_fd_sc_hd__or2_1 _11886_ (.A(_04591_),
    .B(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__mux4_1 _11887_ (.A0(\rbzero.row_render.texu[5] ),
    .A1(\rbzero.row_render.texu[4] ),
    .A2(\rbzero.row_render.texu[3] ),
    .A3(\rbzero.row_render.texu[2] ),
    .S0(_03288_),
    .S1(_04592_),
    .X(_04600_));
 sky130_fd_sc_hd__or2b_1 _11888_ (.A(_04600_),
    .B_N(_04591_),
    .X(_04601_));
 sky130_fd_sc_hd__a31o_1 _11889_ (.A1(_04080_),
    .A2(_04599_),
    .A3(_04601_),
    .B1(_04078_),
    .X(_04602_));
 sky130_fd_sc_hd__or2b_1 _11890_ (.A(\rbzero.row_render.texu[0] ),
    .B_N(_03289_),
    .X(_04603_));
 sky130_fd_sc_hd__nor2_1 _11891_ (.A(_04591_),
    .B(_04592_),
    .Y(_04604_));
 sky130_fd_sc_hd__or2_1 _11892_ (.A(\rbzero.row_render.texu[1] ),
    .B(_03289_),
    .X(_04605_));
 sky130_fd_sc_hd__a31o_1 _11893_ (.A1(_04603_),
    .A2(_04604_),
    .A3(_04605_),
    .B1(_04080_),
    .X(_04606_));
 sky130_fd_sc_hd__nor2_1 _11894_ (.A(_03289_),
    .B(_04604_),
    .Y(_04607_));
 sky130_fd_sc_hd__a21bo_1 _11895_ (.A1(_03289_),
    .A2(_04604_),
    .B1_N(_03782_),
    .X(_04608_));
 sky130_fd_sc_hd__a211o_1 _11896_ (.A1(_04591_),
    .A2(_04592_),
    .B1(_04607_),
    .C1(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__and4b_4 _11897_ (.A_N(o_tex_oeb0),
    .B(_04602_),
    .C(_04606_),
    .D(_04609_),
    .X(_04610_));
 sky130_fd_sc_hd__buf_2 _11898_ (.A(_04610_),
    .X(o_tex_out0));
 sky130_fd_sc_hd__inv_2 _11899_ (.A(net73),
    .Y(o_tex_sclk));
 sky130_fd_sc_hd__clkbuf_2 _11900_ (.A(net9),
    .X(_04611_));
 sky130_fd_sc_hd__or2_1 _11901_ (.A(_04611_),
    .B(o_rgb[14]),
    .X(_04612_));
 sky130_fd_sc_hd__nand2_1 _11902_ (.A(_04611_),
    .B(_04447_),
    .Y(_04613_));
 sky130_fd_sc_hd__a31o_1 _11903_ (.A1(net13),
    .A2(_04612_),
    .A3(_04613_),
    .B1(net12),
    .X(_04614_));
 sky130_fd_sc_hd__nand2_1 _11904_ (.A(net12),
    .B(net13),
    .Y(_04615_));
 sky130_fd_sc_hd__nor2_1 _11905_ (.A(_04611_),
    .B(_04519_),
    .Y(_04616_));
 sky130_fd_sc_hd__a211o_1 _11906_ (.A1(_04611_),
    .A2(o_rgb[23]),
    .B1(_04615_),
    .C1(_04616_),
    .X(_04617_));
 sky130_fd_sc_hd__buf_2 _11907_ (.A(net10),
    .X(_04618_));
 sky130_fd_sc_hd__nor2_1 _11908_ (.A(_04611_),
    .B(_04118_),
    .Y(_04619_));
 sky130_fd_sc_hd__a211o_1 _11909_ (.A1(_04611_),
    .A2(o_rgb[7]),
    .B1(_04619_),
    .C1(net13),
    .X(_04620_));
 sky130_fd_sc_hd__and3_1 _11910_ (.A(_04618_),
    .B(net11),
    .C(_04620_),
    .X(_04621_));
 sky130_fd_sc_hd__and4b_1 _11911_ (.A_N(net14),
    .B(_04614_),
    .C(_04617_),
    .D(_04621_),
    .X(_04622_));
 sky130_fd_sc_hd__nor2_1 _11912_ (.A(net12),
    .B(net11),
    .Y(_04623_));
 sky130_fd_sc_hd__a21o_1 _11913_ (.A1(net10),
    .A2(net11),
    .B1(net12),
    .X(_04624_));
 sky130_fd_sc_hd__and3_1 _11914_ (.A(net14),
    .B(net13),
    .C(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__mux4_1 _11915_ (.A0(_04078_),
    .A1(_03781_),
    .A2(_03784_),
    .A3(_03291_),
    .S0(net9),
    .S1(_04618_),
    .X(_04626_));
 sky130_fd_sc_hd__or2_1 _11916_ (.A(_04625_),
    .B(_04626_),
    .X(_04627_));
 sky130_fd_sc_hd__buf_2 _11917_ (.A(\gpout0.vpos[2] ),
    .X(_04628_));
 sky130_fd_sc_hd__mux4_1 _11918_ (.A0(\gpout0.hpos[2] ),
    .A1(_04080_),
    .A2(_04628_),
    .A3(_04101_),
    .S0(net9),
    .S1(_04625_),
    .X(_04629_));
 sky130_fd_sc_hd__inv_2 _11919_ (.A(net12),
    .Y(_04630_));
 sky130_fd_sc_hd__buf_2 _11920_ (.A(\gpout0.vpos[0] ),
    .X(_04631_));
 sky130_fd_sc_hd__buf_2 _11921_ (.A(\gpout0.vpos[1] ),
    .X(_04632_));
 sky130_fd_sc_hd__mux4_1 _11922_ (.A0(_03288_),
    .A1(_04592_),
    .A2(_04631_),
    .A3(_04632_),
    .S0(net9),
    .S1(_04625_),
    .X(_04633_));
 sky130_fd_sc_hd__o21ba_1 _11923_ (.A1(_04630_),
    .A2(_04633_),
    .B1_N(_04618_),
    .X(_04634_));
 sky130_fd_sc_hd__mux4_1 _11924_ (.A0(_03294_),
    .A1(_03295_),
    .A2(\gpout0.vpos[8] ),
    .A3(_04110_),
    .S0(net9),
    .S1(_04625_),
    .X(_04635_));
 sky130_fd_sc_hd__or2_1 _11925_ (.A(net12),
    .B(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__a32o_1 _11926_ (.A1(_04618_),
    .A2(net12),
    .A3(_04629_),
    .B1(_04634_),
    .B2(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__a22o_1 _11927_ (.A1(_04623_),
    .A2(_04627_),
    .B1(_04637_),
    .B2(net11),
    .X(_04638_));
 sky130_fd_sc_hd__nor2_1 _11928_ (.A(_04630_),
    .B(net11),
    .Y(_04639_));
 sky130_fd_sc_hd__nand2_1 _11929_ (.A(net14),
    .B(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__o22a_1 _11930_ (.A1(net12),
    .A2(net13),
    .B1(_04639_),
    .B2(net14),
    .X(_04641_));
 sky130_fd_sc_hd__and4_1 _11931_ (.A(_04615_),
    .B(_04638_),
    .C(_04640_),
    .D(_04641_),
    .X(_04642_));
 sky130_fd_sc_hd__and2b_1 _11932_ (.A_N(net10),
    .B(net9),
    .X(_04643_));
 sky130_fd_sc_hd__and2b_1 _11933_ (.A_N(net9),
    .B(net10),
    .X(_04644_));
 sky130_fd_sc_hd__and3_1 _11934_ (.A(net48),
    .B(_04611_),
    .C(_04618_),
    .X(_04645_));
 sky130_fd_sc_hd__a221o_1 _11935_ (.A1(o_tex_oeb0),
    .A2(_04643_),
    .B1(_04644_),
    .B2(net47),
    .C1(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__mux4_1 _11936_ (.A0(net42),
    .A1(net44),
    .A2(net43),
    .A3(_04116_),
    .S0(net9),
    .S1(_04618_),
    .X(_04647_));
 sky130_fd_sc_hd__mux4_1 _11937_ (.A0(net49),
    .A1(net40),
    .A2(net39),
    .A3(net41),
    .S0(_04618_),
    .S1(_04611_),
    .X(_04648_));
 sky130_fd_sc_hd__a22o_1 _11938_ (.A1(_04623_),
    .A2(_04647_),
    .B1(_04648_),
    .B2(_04639_),
    .X(_04649_));
 sky130_fd_sc_hd__a31o_1 _11939_ (.A1(_04630_),
    .A2(net11),
    .A3(_04646_),
    .B1(_04649_),
    .X(_04650_));
 sky130_fd_sc_hd__and2b_1 _11940_ (.A_N(net13),
    .B(net14),
    .X(_04651_));
 sky130_fd_sc_hd__nor2_1 _11941_ (.A(_04611_),
    .B(_04618_),
    .Y(_04652_));
 sky130_fd_sc_hd__nor2_1 _11942_ (.A(net14),
    .B(net13),
    .Y(_04653_));
 sky130_fd_sc_hd__a22o_1 _11943_ (.A1(_04115_),
    .A2(_04651_),
    .B1(_04653_),
    .B2(\gpout1.clk_div[1] ),
    .X(_04654_));
 sky130_fd_sc_hd__and3_1 _11944_ (.A(net9),
    .B(_04618_),
    .C(net52),
    .X(_04655_));
 sky130_fd_sc_hd__a221o_1 _11945_ (.A1(net51),
    .A2(_04643_),
    .B1(_04644_),
    .B2(net53),
    .C1(_04655_),
    .X(_04656_));
 sky130_fd_sc_hd__a22o_1 _11946_ (.A1(_04652_),
    .A2(_04654_),
    .B1(_04656_),
    .B2(_04653_),
    .X(_04657_));
 sky130_fd_sc_hd__nand2_1 _11947_ (.A(_04623_),
    .B(_04653_),
    .Y(_04658_));
 sky130_fd_sc_hd__and3b_1 _11948_ (.A_N(\gpout1.clk_div[0] ),
    .B(_04611_),
    .C(_04618_),
    .X(_04659_));
 sky130_fd_sc_hd__a211oi_1 _11949_ (.A1(o_tex_sclk),
    .A2(_04644_),
    .B1(_04658_),
    .C1(_04659_),
    .Y(_04660_));
 sky130_fd_sc_hd__a31o_1 _11950_ (.A1(_04630_),
    .A2(net11),
    .A3(_04657_),
    .B1(_04660_),
    .X(_04661_));
 sky130_fd_sc_hd__a21o_1 _11951_ (.A1(_04650_),
    .A2(_04651_),
    .B1(_04661_),
    .X(_04662_));
 sky130_fd_sc_hd__or3b_1 _11952_ (.A(_04658_),
    .B(o_rgb[15]),
    .C_N(_04652_),
    .X(_04663_));
 sky130_fd_sc_hd__o31a_4 _11953_ (.A1(_04622_),
    .A2(_04642_),
    .A3(_04662_),
    .B1(_04663_),
    .X(o_gpout[1]));
 sky130_fd_sc_hd__buf_2 _11954_ (.A(net16),
    .X(_04664_));
 sky130_fd_sc_hd__buf_2 _11955_ (.A(net15),
    .X(_04665_));
 sky130_fd_sc_hd__nor2_1 _11956_ (.A(net17),
    .B(net18),
    .Y(_04666_));
 sky130_fd_sc_hd__nor2_1 _11957_ (.A(net20),
    .B(net19),
    .Y(_04667_));
 sky130_fd_sc_hd__nand2_1 _11958_ (.A(_04666_),
    .B(_04667_),
    .Y(_04668_));
 sky130_fd_sc_hd__or3_1 _11959_ (.A(_04664_),
    .B(_04665_),
    .C(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__a21o_1 _11960_ (.A1(net16),
    .A2(net17),
    .B1(net18),
    .X(_04670_));
 sky130_fd_sc_hd__and3_1 _11961_ (.A(net20),
    .B(net19),
    .C(_04670_),
    .X(_04671_));
 sky130_fd_sc_hd__mux4_1 _11962_ (.A0(_04078_),
    .A1(_03781_),
    .A2(_03784_),
    .A3(_03291_),
    .S0(_04665_),
    .S1(_04664_),
    .X(_04672_));
 sky130_fd_sc_hd__or2_1 _11963_ (.A(_04671_),
    .B(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__mux4_1 _11964_ (.A0(_04591_),
    .A1(_04080_),
    .A2(_04628_),
    .A3(_04101_),
    .S0(_04665_),
    .S1(_04671_),
    .X(_04674_));
 sky130_fd_sc_hd__mux4_1 _11965_ (.A0(_03294_),
    .A1(_03295_),
    .A2(\gpout0.vpos[8] ),
    .A3(_04110_),
    .S0(net15),
    .S1(_04671_),
    .X(_04675_));
 sky130_fd_sc_hd__o21ba_1 _11966_ (.A1(net18),
    .A2(_04675_),
    .B1_N(_04664_),
    .X(_04676_));
 sky130_fd_sc_hd__inv_2 _11967_ (.A(net18),
    .Y(_04677_));
 sky130_fd_sc_hd__mux4_1 _11968_ (.A0(_03288_),
    .A1(_04592_),
    .A2(_04631_),
    .A3(_04632_),
    .S0(net15),
    .S1(_04671_),
    .X(_04678_));
 sky130_fd_sc_hd__or2_1 _11969_ (.A(_04677_),
    .B(_04678_),
    .X(_04679_));
 sky130_fd_sc_hd__a32o_1 _11970_ (.A1(_04664_),
    .A2(net18),
    .A3(_04674_),
    .B1(_04676_),
    .B2(_04679_),
    .X(_04680_));
 sky130_fd_sc_hd__a22o_1 _11971_ (.A1(_04666_),
    .A2(_04673_),
    .B1(_04680_),
    .B2(net17),
    .X(_04681_));
 sky130_fd_sc_hd__nor2_1 _11972_ (.A(net17),
    .B(_04677_),
    .Y(_04682_));
 sky130_fd_sc_hd__a22oi_1 _11973_ (.A1(net18),
    .A2(net19),
    .B1(_04682_),
    .B2(net20),
    .Y(_04683_));
 sky130_fd_sc_hd__o22a_1 _11974_ (.A1(net18),
    .A2(net19),
    .B1(_04682_),
    .B2(net20),
    .X(_04684_));
 sky130_fd_sc_hd__and3_1 _11975_ (.A(_04681_),
    .B(_04683_),
    .C(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__nand2_1 _11976_ (.A(_04665_),
    .B(_04447_),
    .Y(_04686_));
 sky130_fd_sc_hd__or2_1 _11977_ (.A(_04665_),
    .B(o_rgb[14]),
    .X(_04687_));
 sky130_fd_sc_hd__a31o_1 _11978_ (.A1(net19),
    .A2(_04686_),
    .A3(_04687_),
    .B1(net18),
    .X(_04688_));
 sky130_fd_sc_hd__nor2_1 _11979_ (.A(_04665_),
    .B(_04118_),
    .Y(_04689_));
 sky130_fd_sc_hd__a211o_1 _11980_ (.A1(_04665_),
    .A2(o_rgb[7]),
    .B1(_04689_),
    .C1(net19),
    .X(_04690_));
 sky130_fd_sc_hd__nand2_1 _11981_ (.A(_04665_),
    .B(o_rgb[23]),
    .Y(_04691_));
 sky130_fd_sc_hd__o2111a_1 _11982_ (.A1(_04665_),
    .A2(_04519_),
    .B1(_04691_),
    .C1(net18),
    .D1(net19),
    .X(_04692_));
 sky130_fd_sc_hd__and4bb_1 _11983_ (.A_N(net20),
    .B_N(_04692_),
    .C(_04664_),
    .D(net17),
    .X(_04693_));
 sky130_fd_sc_hd__nor2_1 _11984_ (.A(net16),
    .B(net15),
    .Y(_04694_));
 sky130_fd_sc_hd__and2b_1 _11985_ (.A_N(net19),
    .B(net20),
    .X(_04695_));
 sky130_fd_sc_hd__a22o_1 _11986_ (.A1(\gpout2.clk_div[1] ),
    .A2(_04667_),
    .B1(_04695_),
    .B2(_04115_),
    .X(_04696_));
 sky130_fd_sc_hd__and2b_1 _11987_ (.A_N(net16),
    .B(net15),
    .X(_04697_));
 sky130_fd_sc_hd__and2b_1 _11988_ (.A_N(net15),
    .B(net16),
    .X(_04698_));
 sky130_fd_sc_hd__and3_1 _11989_ (.A(net52),
    .B(_04664_),
    .C(_04665_),
    .X(_04699_));
 sky130_fd_sc_hd__a221o_1 _11990_ (.A1(net51),
    .A2(_04697_),
    .B1(_04698_),
    .B2(net53),
    .C1(_04699_),
    .X(_04700_));
 sky130_fd_sc_hd__a22o_1 _11991_ (.A1(_04694_),
    .A2(_04696_),
    .B1(_04700_),
    .B2(_04667_),
    .X(_04701_));
 sky130_fd_sc_hd__buf_4 _11992_ (.A(net107),
    .X(_04702_));
 sky130_fd_sc_hd__and3_1 _11993_ (.A(\gpout2.clk_div[0] ),
    .B(_04664_),
    .C(net15),
    .X(_04703_));
 sky130_fd_sc_hd__a221o_1 _11994_ (.A1(net45),
    .A2(_04697_),
    .B1(_04698_),
    .B2(_04702_),
    .C1(_04703_),
    .X(_04704_));
 sky130_fd_sc_hd__nor2_1 _11995_ (.A(_04694_),
    .B(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__and3_1 _11996_ (.A(net48),
    .B(_04664_),
    .C(net15),
    .X(_04706_));
 sky130_fd_sc_hd__a221o_1 _11997_ (.A1(o_tex_oeb0),
    .A2(_04697_),
    .B1(_04698_),
    .B2(net47),
    .C1(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__and3_1 _11998_ (.A(_04664_),
    .B(net15),
    .C(_04116_),
    .X(_04708_));
 sky130_fd_sc_hd__a22o_1 _11999_ (.A1(net42),
    .A2(_04694_),
    .B1(_04697_),
    .B2(net44),
    .X(_04709_));
 sky130_fd_sc_hd__a211o_1 _12000_ (.A1(net43),
    .A2(_04698_),
    .B1(_04708_),
    .C1(_04709_),
    .X(_04710_));
 sky130_fd_sc_hd__mux4_1 _12001_ (.A0(net49),
    .A1(net40),
    .A2(net39),
    .A3(net41),
    .S0(_04664_),
    .S1(net15),
    .X(_04711_));
 sky130_fd_sc_hd__a22o_1 _12002_ (.A1(_04666_),
    .A2(_04710_),
    .B1(_04711_),
    .B2(_04682_),
    .X(_04712_));
 sky130_fd_sc_hd__a31o_1 _12003_ (.A1(net17),
    .A2(_04677_),
    .A3(_04707_),
    .B1(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__a2bb2o_1 _12004_ (.A1_N(_04668_),
    .A2_N(_04705_),
    .B1(_04695_),
    .B2(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__a31o_1 _12005_ (.A1(net17),
    .A2(_04677_),
    .A3(_04701_),
    .B1(_04714_),
    .X(_04715_));
 sky130_fd_sc_hd__a31o_1 _12006_ (.A1(_04688_),
    .A2(_04690_),
    .A3(_04693_),
    .B1(_04715_),
    .X(_04716_));
 sky130_fd_sc_hd__o22a_2 _12007_ (.A1(o_rgb[6]),
    .A2(_04669_),
    .B1(_04685_),
    .B2(_04716_),
    .X(o_gpout[2]));
 sky130_fd_sc_hd__buf_2 _12008_ (.A(net3),
    .X(_04717_));
 sky130_fd_sc_hd__buf_2 _12009_ (.A(net4),
    .X(_04718_));
 sky130_fd_sc_hd__nor2_1 _12010_ (.A(net5),
    .B(net6),
    .Y(_04719_));
 sky130_fd_sc_hd__nor2_1 _12011_ (.A(net8),
    .B(net7),
    .Y(_04720_));
 sky130_fd_sc_hd__nand2_1 _12012_ (.A(_04719_),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__nand2_1 _12013_ (.A(_04717_),
    .B(_04447_),
    .Y(_04722_));
 sky130_fd_sc_hd__o211a_1 _12014_ (.A1(_04717_),
    .A2(o_rgb[14]),
    .B1(_04722_),
    .C1(net7),
    .X(_04723_));
 sky130_fd_sc_hd__nor2_1 _12015_ (.A(_04717_),
    .B(_04118_),
    .Y(_04724_));
 sky130_fd_sc_hd__a211o_1 _12016_ (.A1(_04717_),
    .A2(o_rgb[7]),
    .B1(_04724_),
    .C1(net7),
    .X(_04725_));
 sky130_fd_sc_hd__nand2_1 _12017_ (.A(_04717_),
    .B(o_rgb[23]),
    .Y(_04726_));
 sky130_fd_sc_hd__o2111a_1 _12018_ (.A1(_04717_),
    .A2(_04519_),
    .B1(_04726_),
    .C1(net6),
    .D1(net7),
    .X(_04727_));
 sky130_fd_sc_hd__and4bb_1 _12019_ (.A_N(net8),
    .B_N(_04727_),
    .C(_04718_),
    .D(net5),
    .X(_04728_));
 sky130_fd_sc_hd__o211a_1 _12020_ (.A1(net6),
    .A2(_04723_),
    .B1(_04725_),
    .C1(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__a21o_1 _12021_ (.A1(net4),
    .A2(net5),
    .B1(net6),
    .X(_04730_));
 sky130_fd_sc_hd__and3_1 _12022_ (.A(net8),
    .B(net7),
    .C(_04730_),
    .X(_04731_));
 sky130_fd_sc_hd__mux4_1 _12023_ (.A0(\gpout0.hpos[2] ),
    .A1(_04080_),
    .A2(_04628_),
    .A3(_04101_),
    .S0(net3),
    .S1(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__mux4_1 _12024_ (.A0(_03294_),
    .A1(_03295_),
    .A2(\gpout0.vpos[8] ),
    .A3(_04110_),
    .S0(net3),
    .S1(_04731_),
    .X(_04733_));
 sky130_fd_sc_hd__o21ba_1 _12025_ (.A1(net6),
    .A2(_04733_),
    .B1_N(_04718_),
    .X(_04734_));
 sky130_fd_sc_hd__inv_2 _12026_ (.A(net6),
    .Y(_04735_));
 sky130_fd_sc_hd__mux4_1 _12027_ (.A0(_03288_),
    .A1(\gpout0.hpos[1] ),
    .A2(\gpout0.vpos[0] ),
    .A3(_04632_),
    .S0(net3),
    .S1(_04731_),
    .X(_04736_));
 sky130_fd_sc_hd__or2_1 _12028_ (.A(_04735_),
    .B(_04736_),
    .X(_04737_));
 sky130_fd_sc_hd__a32o_1 _12029_ (.A1(_04718_),
    .A2(net6),
    .A3(_04732_),
    .B1(_04734_),
    .B2(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__mux4_1 _12030_ (.A0(_04078_),
    .A1(_03781_),
    .A2(_04106_),
    .A3(_04104_),
    .S0(_04717_),
    .S1(_04731_),
    .X(_04739_));
 sky130_fd_sc_hd__mux4_1 _12031_ (.A0(_03784_),
    .A1(_03291_),
    .A2(\gpout0.vpos[6] ),
    .A3(\gpout0.vpos[7] ),
    .S0(net3),
    .S1(_04731_),
    .X(_04740_));
 sky130_fd_sc_hd__mux2_1 _12032_ (.A0(_04739_),
    .A1(_04740_),
    .S(_04718_),
    .X(_04741_));
 sky130_fd_sc_hd__a22o_1 _12033_ (.A1(net5),
    .A2(_04738_),
    .B1(_04719_),
    .B2(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__nor2_1 _12034_ (.A(net5),
    .B(_04735_),
    .Y(_04743_));
 sky130_fd_sc_hd__a22oi_1 _12035_ (.A1(net6),
    .A2(net7),
    .B1(_04743_),
    .B2(net8),
    .Y(_04744_));
 sky130_fd_sc_hd__o22a_1 _12036_ (.A1(net6),
    .A2(net7),
    .B1(_04743_),
    .B2(net8),
    .X(_04745_));
 sky130_fd_sc_hd__and3_1 _12037_ (.A(_04742_),
    .B(_04744_),
    .C(_04745_),
    .X(_04746_));
 sky130_fd_sc_hd__nor2_1 _12038_ (.A(_04718_),
    .B(_03292_),
    .Y(_04747_));
 sky130_fd_sc_hd__and2b_1 _12039_ (.A_N(net3),
    .B(_04718_),
    .X(_04748_));
 sky130_fd_sc_hd__and2_1 _12040_ (.A(net3),
    .B(_04718_),
    .X(_04749_));
 sky130_fd_sc_hd__nor2_1 _12041_ (.A(net3),
    .B(net4),
    .Y(_04750_));
 sky130_fd_sc_hd__a221o_1 _12042_ (.A1(_04702_),
    .A2(_04748_),
    .B1(_04749_),
    .B2(\gpout0.clk_div[0] ),
    .C1(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__o21ba_1 _12043_ (.A1(_04747_),
    .A2(_04751_),
    .B1_N(_04721_),
    .X(_04752_));
 sky130_fd_sc_hd__and2b_1 _12044_ (.A_N(net7),
    .B(net8),
    .X(_04753_));
 sky130_fd_sc_hd__a22o_1 _12045_ (.A1(_04115_),
    .A2(_04753_),
    .B1(_04720_),
    .B2(\gpout0.clk_div[1] ),
    .X(_04754_));
 sky130_fd_sc_hd__and2b_1 _12046_ (.A_N(net4),
    .B(net3),
    .X(_04755_));
 sky130_fd_sc_hd__and3_1 _12047_ (.A(net52),
    .B(_04717_),
    .C(_04718_),
    .X(_04756_));
 sky130_fd_sc_hd__a221o_1 _12048_ (.A1(net53),
    .A2(_04748_),
    .B1(_04755_),
    .B2(net51),
    .C1(_04756_),
    .X(_04757_));
 sky130_fd_sc_hd__a22o_1 _12049_ (.A1(_04750_),
    .A2(_04754_),
    .B1(_04757_),
    .B2(_04720_),
    .X(_04758_));
 sky130_fd_sc_hd__a22o_1 _12050_ (.A1(net47),
    .A2(_04748_),
    .B1(_04749_),
    .B2(net48),
    .X(_04759_));
 sky130_fd_sc_hd__a21o_1 _12051_ (.A1(o_tex_oeb0),
    .A2(_04755_),
    .B1(_04759_),
    .X(_04760_));
 sky130_fd_sc_hd__a22o_1 _12052_ (.A1(net42),
    .A2(_04750_),
    .B1(_04755_),
    .B2(net44),
    .X(_04761_));
 sky130_fd_sc_hd__a221o_1 _12053_ (.A1(net43),
    .A2(_04748_),
    .B1(_04749_),
    .B2(_04116_),
    .C1(_04761_),
    .X(_04762_));
 sky130_fd_sc_hd__mux4_1 _12054_ (.A0(net49),
    .A1(net40),
    .A2(net39),
    .A3(net41),
    .S0(_04718_),
    .S1(_04717_),
    .X(_04763_));
 sky130_fd_sc_hd__a22o_1 _12055_ (.A1(_04719_),
    .A2(_04762_),
    .B1(_04763_),
    .B2(_04743_),
    .X(_04764_));
 sky130_fd_sc_hd__a31o_1 _12056_ (.A1(net5),
    .A2(_04735_),
    .A3(_04760_),
    .B1(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__a32o_1 _12057_ (.A1(net5),
    .A2(_04735_),
    .A3(_04758_),
    .B1(_04765_),
    .B2(_04753_),
    .X(_04766_));
 sky130_fd_sc_hd__or4_1 _12058_ (.A(_04729_),
    .B(_04746_),
    .C(_04752_),
    .D(_04766_),
    .X(_04767_));
 sky130_fd_sc_hd__o41a_4 _12059_ (.A1(_04717_),
    .A2(_04718_),
    .A3(o_rgb[14]),
    .A4(_04721_),
    .B1(_04767_),
    .X(o_gpout[0]));
 sky130_fd_sc_hd__buf_2 _12060_ (.A(net21),
    .X(_04768_));
 sky130_fd_sc_hd__nand2_1 _12061_ (.A(_04768_),
    .B(_04447_),
    .Y(_04769_));
 sky130_fd_sc_hd__o211a_1 _12062_ (.A1(_04768_),
    .A2(o_rgb[14]),
    .B1(_04769_),
    .C1(net25),
    .X(_04770_));
 sky130_fd_sc_hd__nor2_1 _12063_ (.A(_04768_),
    .B(_04118_),
    .Y(_04771_));
 sky130_fd_sc_hd__a211o_1 _12064_ (.A1(_04768_),
    .A2(o_rgb[7]),
    .B1(_04771_),
    .C1(net25),
    .X(_04772_));
 sky130_fd_sc_hd__buf_2 _12065_ (.A(net22),
    .X(_04773_));
 sky130_fd_sc_hd__and4b_1 _12066_ (.A_N(net26),
    .B(_04772_),
    .C(_04773_),
    .D(net23),
    .X(_04774_));
 sky130_fd_sc_hd__nand2_1 _12067_ (.A(net24),
    .B(net25),
    .Y(_04775_));
 sky130_fd_sc_hd__nor2_1 _12068_ (.A(_04768_),
    .B(_04519_),
    .Y(_04776_));
 sky130_fd_sc_hd__a211o_1 _12069_ (.A1(_04768_),
    .A2(o_rgb[23]),
    .B1(_04775_),
    .C1(_04776_),
    .X(_04777_));
 sky130_fd_sc_hd__o211a_1 _12070_ (.A1(net24),
    .A2(_04770_),
    .B1(_04774_),
    .C1(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__nor2_1 _12071_ (.A(net24),
    .B(net23),
    .Y(_04779_));
 sky130_fd_sc_hd__a21o_1 _12072_ (.A1(net22),
    .A2(net23),
    .B1(net24),
    .X(_04780_));
 sky130_fd_sc_hd__and3_1 _12073_ (.A(net26),
    .B(net25),
    .C(_04780_),
    .X(_04781_));
 sky130_fd_sc_hd__mux4_1 _12074_ (.A0(_04078_),
    .A1(_03781_),
    .A2(_03784_),
    .A3(_03291_),
    .S0(net21),
    .S1(_04773_),
    .X(_04782_));
 sky130_fd_sc_hd__or2_1 _12075_ (.A(_04781_),
    .B(_04782_),
    .X(_04783_));
 sky130_fd_sc_hd__mux4_1 _12076_ (.A0(_04591_),
    .A1(_04080_),
    .A2(_04628_),
    .A3(_04101_),
    .S0(net21),
    .S1(_04781_),
    .X(_04784_));
 sky130_fd_sc_hd__inv_2 _12077_ (.A(net24),
    .Y(_04785_));
 sky130_fd_sc_hd__mux4_1 _12078_ (.A0(_03288_),
    .A1(\gpout0.hpos[1] ),
    .A2(_04631_),
    .A3(_04632_),
    .S0(net21),
    .S1(_04781_),
    .X(_04786_));
 sky130_fd_sc_hd__mux4_1 _12079_ (.A0(_03294_),
    .A1(_03295_),
    .A2(\gpout0.vpos[8] ),
    .A3(_04110_),
    .S0(net21),
    .S1(_04781_),
    .X(_04787_));
 sky130_fd_sc_hd__or2_1 _12080_ (.A(net24),
    .B(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__inv_2 _12081_ (.A(_04773_),
    .Y(_04789_));
 sky130_fd_sc_hd__o211a_1 _12082_ (.A1(_04785_),
    .A2(_04786_),
    .B1(_04788_),
    .C1(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__a31o_1 _12083_ (.A1(_04773_),
    .A2(net24),
    .A3(_04784_),
    .B1(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__a22o_1 _12084_ (.A1(_04779_),
    .A2(_04783_),
    .B1(_04791_),
    .B2(net23),
    .X(_04792_));
 sky130_fd_sc_hd__nor2_1 _12085_ (.A(_04785_),
    .B(net23),
    .Y(_04793_));
 sky130_fd_sc_hd__nand2_1 _12086_ (.A(net26),
    .B(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__o22a_1 _12087_ (.A1(net24),
    .A2(net25),
    .B1(_04793_),
    .B2(net26),
    .X(_04795_));
 sky130_fd_sc_hd__and4_1 _12088_ (.A(_04775_),
    .B(_04792_),
    .C(_04794_),
    .D(_04795_),
    .X(_04796_));
 sky130_fd_sc_hd__and2b_1 _12089_ (.A_N(net25),
    .B(net26),
    .X(_04797_));
 sky130_fd_sc_hd__and2_1 _12090_ (.A(_04789_),
    .B(net21),
    .X(_04798_));
 sky130_fd_sc_hd__nor2_1 _12091_ (.A(_04789_),
    .B(_04768_),
    .Y(_04799_));
 sky130_fd_sc_hd__and3_1 _12092_ (.A(net48),
    .B(_04773_),
    .C(_04768_),
    .X(_04800_));
 sky130_fd_sc_hd__a221o_1 _12093_ (.A1(o_tex_oeb0),
    .A2(_04798_),
    .B1(_04799_),
    .B2(net47),
    .C1(_04800_),
    .X(_04801_));
 sky130_fd_sc_hd__and3_1 _12094_ (.A(_04773_),
    .B(net21),
    .C(_04116_),
    .X(_04802_));
 sky130_fd_sc_hd__nor2_1 _12095_ (.A(_04773_),
    .B(net21),
    .Y(_04803_));
 sky130_fd_sc_hd__a22o_1 _12096_ (.A1(net44),
    .A2(_04798_),
    .B1(_04803_),
    .B2(net42),
    .X(_04804_));
 sky130_fd_sc_hd__a211o_1 _12097_ (.A1(net43),
    .A2(_04799_),
    .B1(_04802_),
    .C1(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__mux4_1 _12098_ (.A0(net49),
    .A1(net40),
    .A2(net39),
    .A3(net41),
    .S0(_04773_),
    .S1(_04768_),
    .X(_04806_));
 sky130_fd_sc_hd__a22o_1 _12099_ (.A1(_04779_),
    .A2(_04805_),
    .B1(_04806_),
    .B2(_04793_),
    .X(_04807_));
 sky130_fd_sc_hd__a31o_1 _12100_ (.A1(_04785_),
    .A2(net23),
    .A3(_04801_),
    .B1(_04807_),
    .X(_04808_));
 sky130_fd_sc_hd__nor2_1 _12101_ (.A(net26),
    .B(net25),
    .Y(_04809_));
 sky130_fd_sc_hd__a22o_1 _12102_ (.A1(_04115_),
    .A2(_04797_),
    .B1(_04809_),
    .B2(\gpout3.clk_div[1] ),
    .X(_04810_));
 sky130_fd_sc_hd__and3_1 _12103_ (.A(net52),
    .B(_04773_),
    .C(_04768_),
    .X(_04811_));
 sky130_fd_sc_hd__a221o_1 _12104_ (.A1(net51),
    .A2(_04798_),
    .B1(_04799_),
    .B2(net53),
    .C1(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__a22o_1 _12105_ (.A1(_04803_),
    .A2(_04810_),
    .B1(_04812_),
    .B2(_04809_),
    .X(_04813_));
 sky130_fd_sc_hd__and3_1 _12106_ (.A(_04773_),
    .B(net21),
    .C(\gpout3.clk_div[0] ),
    .X(_04814_));
 sky130_fd_sc_hd__a221o_1 _12107_ (.A1(net46),
    .A2(_04798_),
    .B1(_04799_),
    .B2(_04702_),
    .C1(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__o211a_1 _12108_ (.A1(_04803_),
    .A2(_04815_),
    .B1(_04809_),
    .C1(_04779_),
    .X(_04816_));
 sky130_fd_sc_hd__a31o_1 _12109_ (.A1(_04785_),
    .A2(net23),
    .A3(_04813_),
    .B1(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__a21o_1 _12110_ (.A1(_04797_),
    .A2(_04808_),
    .B1(_04817_),
    .X(_04818_));
 sky130_fd_sc_hd__nand4b_1 _12111_ (.A_N(o_rgb[7]),
    .B(_04779_),
    .C(_04803_),
    .D(_04809_),
    .Y(_04819_));
 sky130_fd_sc_hd__o31a_4 _12112_ (.A1(_04778_),
    .A2(_04796_),
    .A3(_04818_),
    .B1(_04819_),
    .X(o_gpout[3]));
 sky130_fd_sc_hd__buf_2 _12113_ (.A(net27),
    .X(_04820_));
 sky130_fd_sc_hd__nand2_1 _12114_ (.A(_04820_),
    .B(_04447_),
    .Y(_04821_));
 sky130_fd_sc_hd__o211a_1 _12115_ (.A1(_04820_),
    .A2(o_rgb[14]),
    .B1(_04821_),
    .C1(net31),
    .X(_04822_));
 sky130_fd_sc_hd__nor2_1 _12116_ (.A(_04820_),
    .B(_04118_),
    .Y(_04823_));
 sky130_fd_sc_hd__a211o_1 _12117_ (.A1(_04820_),
    .A2(o_rgb[7]),
    .B1(_04823_),
    .C1(net31),
    .X(_04824_));
 sky130_fd_sc_hd__buf_2 _12118_ (.A(net28),
    .X(_04825_));
 sky130_fd_sc_hd__and4b_1 _12119_ (.A_N(net32),
    .B(_04824_),
    .C(_04825_),
    .D(net29),
    .X(_04826_));
 sky130_fd_sc_hd__o211a_1 _12120_ (.A1(_04820_),
    .A2(_04519_),
    .B1(net31),
    .C1(net30),
    .X(_04827_));
 sky130_fd_sc_hd__a21bo_1 _12121_ (.A1(_04820_),
    .A2(o_rgb[23]),
    .B1_N(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__o211a_1 _12122_ (.A1(net30),
    .A2(_04822_),
    .B1(_04826_),
    .C1(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__nor2_1 _12123_ (.A(net30),
    .B(net29),
    .Y(_04830_));
 sky130_fd_sc_hd__a21o_1 _12124_ (.A1(net28),
    .A2(net29),
    .B1(net30),
    .X(_04831_));
 sky130_fd_sc_hd__and3_1 _12125_ (.A(net32),
    .B(net31),
    .C(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__mux4_1 _12126_ (.A0(_04078_),
    .A1(_03781_),
    .A2(_03784_),
    .A3(_03291_),
    .S0(net27),
    .S1(_04825_),
    .X(_04833_));
 sky130_fd_sc_hd__or2_1 _12127_ (.A(_04832_),
    .B(_04833_),
    .X(_04834_));
 sky130_fd_sc_hd__mux4_1 _12128_ (.A0(_04591_),
    .A1(_04080_),
    .A2(_04628_),
    .A3(_04101_),
    .S0(_04820_),
    .S1(_04832_),
    .X(_04835_));
 sky130_fd_sc_hd__inv_2 _12129_ (.A(net30),
    .Y(_04836_));
 sky130_fd_sc_hd__mux4_1 _12130_ (.A0(_03288_),
    .A1(\gpout0.hpos[1] ),
    .A2(_04631_),
    .A3(_04632_),
    .S0(net27),
    .S1(_04832_),
    .X(_04837_));
 sky130_fd_sc_hd__mux4_1 _12131_ (.A0(_03294_),
    .A1(_03295_),
    .A2(\gpout0.vpos[8] ),
    .A3(_04110_),
    .S0(net27),
    .S1(_04832_),
    .X(_04838_));
 sky130_fd_sc_hd__or2_1 _12132_ (.A(net30),
    .B(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__inv_2 _12133_ (.A(_04825_),
    .Y(_04840_));
 sky130_fd_sc_hd__o211a_1 _12134_ (.A1(_04836_),
    .A2(_04837_),
    .B1(_04839_),
    .C1(_04840_),
    .X(_04841_));
 sky130_fd_sc_hd__a31o_1 _12135_ (.A1(_04825_),
    .A2(net30),
    .A3(_04835_),
    .B1(_04841_),
    .X(_04842_));
 sky130_fd_sc_hd__a22o_1 _12136_ (.A1(_04830_),
    .A2(_04834_),
    .B1(_04842_),
    .B2(net29),
    .X(_04843_));
 sky130_fd_sc_hd__nor2_1 _12137_ (.A(_04836_),
    .B(net29),
    .Y(_04844_));
 sky130_fd_sc_hd__a22oi_1 _12138_ (.A1(net30),
    .A2(net31),
    .B1(_04844_),
    .B2(net32),
    .Y(_04845_));
 sky130_fd_sc_hd__o22a_1 _12139_ (.A1(net30),
    .A2(net31),
    .B1(_04844_),
    .B2(net32),
    .X(_04846_));
 sky130_fd_sc_hd__and3_1 _12140_ (.A(_04843_),
    .B(_04845_),
    .C(_04846_),
    .X(_04847_));
 sky130_fd_sc_hd__and2_1 _12141_ (.A(_04840_),
    .B(net27),
    .X(_04848_));
 sky130_fd_sc_hd__nor2_1 _12142_ (.A(_04840_),
    .B(_04820_),
    .Y(_04849_));
 sky130_fd_sc_hd__and3_1 _12143_ (.A(net48),
    .B(_04825_),
    .C(_04820_),
    .X(_04850_));
 sky130_fd_sc_hd__a221o_1 _12144_ (.A1(o_tex_oeb0),
    .A2(_04848_),
    .B1(_04849_),
    .B2(net47),
    .C1(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__and3_1 _12145_ (.A(_04825_),
    .B(net27),
    .C(_04116_),
    .X(_04852_));
 sky130_fd_sc_hd__nor2_1 _12146_ (.A(_04825_),
    .B(net27),
    .Y(_04853_));
 sky130_fd_sc_hd__a22o_1 _12147_ (.A1(net44),
    .A2(_04848_),
    .B1(_04853_),
    .B2(net42),
    .X(_04854_));
 sky130_fd_sc_hd__a211o_1 _12148_ (.A1(net43),
    .A2(_04849_),
    .B1(_04852_),
    .C1(_04854_),
    .X(_04855_));
 sky130_fd_sc_hd__mux4_1 _12149_ (.A0(net49),
    .A1(net40),
    .A2(net39),
    .A3(net41),
    .S0(_04825_),
    .S1(_04820_),
    .X(_04856_));
 sky130_fd_sc_hd__a22o_1 _12150_ (.A1(_04830_),
    .A2(_04855_),
    .B1(_04856_),
    .B2(_04844_),
    .X(_04857_));
 sky130_fd_sc_hd__a31o_1 _12151_ (.A1(_04836_),
    .A2(net29),
    .A3(_04851_),
    .B1(_04857_),
    .X(_04858_));
 sky130_fd_sc_hd__and2b_1 _12152_ (.A_N(net31),
    .B(net32),
    .X(_04859_));
 sky130_fd_sc_hd__nor2_1 _12153_ (.A(net32),
    .B(net31),
    .Y(_04860_));
 sky130_fd_sc_hd__a22o_1 _12154_ (.A1(_04115_),
    .A2(_04859_),
    .B1(_04860_),
    .B2(\gpout4.clk_div[1] ),
    .X(_04861_));
 sky130_fd_sc_hd__and3_1 _12155_ (.A(net52),
    .B(_04825_),
    .C(net27),
    .X(_04862_));
 sky130_fd_sc_hd__a221o_1 _12156_ (.A1(net51),
    .A2(_04848_),
    .B1(_04849_),
    .B2(net53),
    .C1(_04862_),
    .X(_04863_));
 sky130_fd_sc_hd__a22o_1 _12157_ (.A1(_04853_),
    .A2(_04861_),
    .B1(_04863_),
    .B2(_04860_),
    .X(_04864_));
 sky130_fd_sc_hd__and3_1 _12158_ (.A(_04825_),
    .B(net27),
    .C(\gpout4.clk_div[0] ),
    .X(_04865_));
 sky130_fd_sc_hd__a221o_1 _12159_ (.A1(net2),
    .A2(_04848_),
    .B1(_04849_),
    .B2(_04702_),
    .C1(_04865_),
    .X(_04866_));
 sky130_fd_sc_hd__o211a_1 _12160_ (.A1(_04853_),
    .A2(_04866_),
    .B1(_04860_),
    .C1(_04830_),
    .X(_04867_));
 sky130_fd_sc_hd__a31o_1 _12161_ (.A1(_04836_),
    .A2(net29),
    .A3(_04864_),
    .B1(_04867_),
    .X(_04868_));
 sky130_fd_sc_hd__a21o_1 _12162_ (.A1(_04858_),
    .A2(_04859_),
    .B1(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__nand3_1 _12163_ (.A(_04830_),
    .B(_04853_),
    .C(_04860_),
    .Y(_04870_));
 sky130_fd_sc_hd__o32a_4 _12164_ (.A1(_04829_),
    .A2(_04847_),
    .A3(_04869_),
    .B1(_04870_),
    .B2(o_rgb[22]),
    .X(o_gpout[4]));
 sky130_fd_sc_hd__inv_2 _12165_ (.A(net36),
    .Y(_04871_));
 sky130_fd_sc_hd__nor2_1 _12166_ (.A(_04871_),
    .B(net35),
    .Y(_04872_));
 sky130_fd_sc_hd__buf_2 _12167_ (.A(net34),
    .X(_04873_));
 sky130_fd_sc_hd__buf_2 _12168_ (.A(net33),
    .X(_04874_));
 sky130_fd_sc_hd__a21o_1 _12169_ (.A1(net34),
    .A2(net35),
    .B1(net36),
    .X(_04875_));
 sky130_fd_sc_hd__and3_1 _12170_ (.A(net38),
    .B(net37),
    .C(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__mux4_1 _12171_ (.A0(_04591_),
    .A1(_04080_),
    .A2(_04628_),
    .A3(_04101_),
    .S0(_04874_),
    .S1(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__mux4_1 _12172_ (.A0(_03294_),
    .A1(_03295_),
    .A2(\gpout0.vpos[8] ),
    .A3(_04110_),
    .S0(_04874_),
    .S1(_04876_),
    .X(_04878_));
 sky130_fd_sc_hd__o21ba_1 _12173_ (.A1(net36),
    .A2(_04878_),
    .B1_N(_04873_),
    .X(_04879_));
 sky130_fd_sc_hd__mux4_1 _12174_ (.A0(_03288_),
    .A1(_04592_),
    .A2(_04631_),
    .A3(_04632_),
    .S0(_04874_),
    .S1(_04876_),
    .X(_04880_));
 sky130_fd_sc_hd__or2_1 _12175_ (.A(_04871_),
    .B(_04880_),
    .X(_04881_));
 sky130_fd_sc_hd__a32o_1 _12176_ (.A1(_04873_),
    .A2(net36),
    .A3(_04877_),
    .B1(_04879_),
    .B2(_04881_),
    .X(_04882_));
 sky130_fd_sc_hd__buf_2 _12177_ (.A(_04874_),
    .X(_04883_));
 sky130_fd_sc_hd__mux4_1 _12178_ (.A0(_04078_),
    .A1(_03781_),
    .A2(_03784_),
    .A3(_03291_),
    .S0(_04883_),
    .S1(_04873_),
    .X(_04884_));
 sky130_fd_sc_hd__nor2_1 _12179_ (.A(net36),
    .B(net35),
    .Y(_04885_));
 sky130_fd_sc_hd__o21a_1 _12180_ (.A1(_04876_),
    .A2(_04884_),
    .B1(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__a21oi_1 _12181_ (.A1(net35),
    .A2(_04882_),
    .B1(_04886_),
    .Y(_04887_));
 sky130_fd_sc_hd__a221oi_1 _12182_ (.A1(net36),
    .A2(net37),
    .B1(_04872_),
    .B2(net38),
    .C1(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__o221a_1 _12183_ (.A1(net36),
    .A2(net37),
    .B1(_04872_),
    .B2(net38),
    .C1(_04888_),
    .X(_04889_));
 sky130_fd_sc_hd__or2_1 _12184_ (.A(_04883_),
    .B(o_rgb[14]),
    .X(_04890_));
 sky130_fd_sc_hd__nand2_1 _12185_ (.A(_04883_),
    .B(_04447_),
    .Y(_04891_));
 sky130_fd_sc_hd__a31o_1 _12186_ (.A1(net37),
    .A2(_04890_),
    .A3(_04891_),
    .B1(net36),
    .X(_04892_));
 sky130_fd_sc_hd__nor2_1 _12187_ (.A(_04883_),
    .B(_04118_),
    .Y(_04893_));
 sky130_fd_sc_hd__a211o_1 _12188_ (.A1(_04883_),
    .A2(o_rgb[7]),
    .B1(_04893_),
    .C1(net37),
    .X(_04894_));
 sky130_fd_sc_hd__inv_2 _12189_ (.A(net38),
    .Y(_04895_));
 sky130_fd_sc_hd__o211a_1 _12190_ (.A1(_04883_),
    .A2(_04519_),
    .B1(net37),
    .C1(net36),
    .X(_04896_));
 sky130_fd_sc_hd__a21bo_1 _12191_ (.A1(_04883_),
    .A2(o_rgb[23]),
    .B1_N(_04896_),
    .X(_04897_));
 sky130_fd_sc_hd__and4_1 _12192_ (.A(_04873_),
    .B(net35),
    .C(_04895_),
    .D(_04897_),
    .X(_04898_));
 sky130_fd_sc_hd__and2b_1 _12193_ (.A_N(net33),
    .B(net34),
    .X(_04899_));
 sky130_fd_sc_hd__and2b_1 _12194_ (.A_N(net34),
    .B(_04874_),
    .X(_04900_));
 sky130_fd_sc_hd__and3_1 _12195_ (.A(net48),
    .B(net34),
    .C(_04874_),
    .X(_04901_));
 sky130_fd_sc_hd__a221o_1 _12196_ (.A1(net47),
    .A2(_04899_),
    .B1(_04900_),
    .B2(o_tex_oeb0),
    .C1(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__mux4_1 _12197_ (.A0(net49),
    .A1(net40),
    .A2(net39),
    .A3(net41),
    .S0(net34),
    .S1(_04874_),
    .X(_04903_));
 sky130_fd_sc_hd__a22o_1 _12198_ (.A1(net43),
    .A2(_04899_),
    .B1(_04900_),
    .B2(net44),
    .X(_04904_));
 sky130_fd_sc_hd__a31o_1 _12199_ (.A1(_04873_),
    .A2(_04874_),
    .A3(_04116_),
    .B1(_04904_),
    .X(_04905_));
 sky130_fd_sc_hd__a221o_1 _12200_ (.A1(_04872_),
    .A2(_04903_),
    .B1(_04905_),
    .B2(_04885_),
    .C1(_04895_),
    .X(_04906_));
 sky130_fd_sc_hd__nand2_1 _12201_ (.A(net35),
    .B(_04115_),
    .Y(_04907_));
 sky130_fd_sc_hd__o2bb2a_1 _12202_ (.A1_N(net42),
    .A2_N(_04885_),
    .B1(_04907_),
    .B2(net36),
    .X(_04908_));
 sky130_fd_sc_hd__nor3_1 _12203_ (.A(_04873_),
    .B(_04883_),
    .C(_04908_),
    .Y(_04909_));
 sky130_fd_sc_hd__a311o_1 _12204_ (.A1(_04871_),
    .A2(net35),
    .A3(_04902_),
    .B1(_04906_),
    .C1(_04909_),
    .X(_04910_));
 sky130_fd_sc_hd__mux4_1 _12205_ (.A0(\gpout5.clk_div[1] ),
    .A1(net51),
    .A2(net53),
    .A3(net52),
    .S0(_04883_),
    .S1(_04873_),
    .X(_04911_));
 sky130_fd_sc_hd__a21oi_1 _12206_ (.A1(o_tex_sclk),
    .A2(_04873_),
    .B1(_04874_),
    .Y(_04912_));
 sky130_fd_sc_hd__a31o_1 _12207_ (.A1(_04873_),
    .A2(_04874_),
    .A3(\gpout5.clk_div[0] ),
    .B1(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__a21o_1 _12208_ (.A1(_04885_),
    .A2(_04913_),
    .B1(net38),
    .X(_04914_));
 sky130_fd_sc_hd__a31o_1 _12209_ (.A1(_04871_),
    .A2(net35),
    .A3(_04911_),
    .B1(_04914_),
    .X(_04915_));
 sky130_fd_sc_hd__and3b_1 _12210_ (.A_N(net37),
    .B(_04910_),
    .C(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__a31o_1 _12211_ (.A1(_04892_),
    .A2(_04894_),
    .A3(_04898_),
    .B1(_04916_),
    .X(_04917_));
 sky130_fd_sc_hd__or4_1 _12212_ (.A(_04873_),
    .B(_04883_),
    .C(net38),
    .D(net37),
    .X(_04918_));
 sky130_fd_sc_hd__or3b_1 _12213_ (.A(_04918_),
    .B(o_rgb[23]),
    .C_N(_04885_),
    .X(_04919_));
 sky130_fd_sc_hd__o21a_2 _12214_ (.A1(_04889_),
    .A2(_04917_),
    .B1(_04919_),
    .X(o_gpout[5]));
 sky130_fd_sc_hd__inv_2 _12215_ (.A(\rbzero.hsync ),
    .Y(o_hsync));
 sky130_fd_sc_hd__buf_4 _12216_ (.A(_03292_),
    .X(_04920_));
 sky130_fd_sc_hd__and3_1 _12217_ (.A(o_vsync),
    .B(\rbzero.wall_tracer.state[12] ),
    .C(_04920_),
    .X(_04921_));
 sky130_fd_sc_hd__clkbuf_1 _12218_ (.A(_04921_),
    .X(_00001_));
 sky130_fd_sc_hd__and3_1 _12219_ (.A(o_vsync),
    .B(\rbzero.wall_tracer.state[2] ),
    .C(_04920_),
    .X(_04922_));
 sky130_fd_sc_hd__clkbuf_1 _12220_ (.A(_04922_),
    .X(_00006_));
 sky130_fd_sc_hd__and3_1 _12221_ (.A(o_vsync),
    .B(\rbzero.wall_tracer.state[7] ),
    .C(_04920_),
    .X(_04923_));
 sky130_fd_sc_hd__clkbuf_1 _12222_ (.A(_04923_),
    .X(_00002_));
 sky130_fd_sc_hd__nor2_1 _12223_ (.A(_03791_),
    .B(_03730_),
    .Y(_00003_));
 sky130_fd_sc_hd__and3_1 _12224_ (.A(o_vsync),
    .B(\rbzero.wall_tracer.state[9] ),
    .C(_03292_),
    .X(_04924_));
 sky130_fd_sc_hd__clkbuf_4 _12225_ (.A(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__buf_4 _12226_ (.A(_04925_),
    .X(_00004_));
 sky130_fd_sc_hd__nor2_1 _12227_ (.A(_03817_),
    .B(_03730_),
    .Y(_00005_));
 sky130_fd_sc_hd__and3_1 _12228_ (.A(o_vsync),
    .B(\rbzero.wall_tracer.state[5] ),
    .C(_04920_),
    .X(_04926_));
 sky130_fd_sc_hd__clkbuf_1 _12229_ (.A(_04926_),
    .X(_00009_));
 sky130_fd_sc_hd__inv_2 _12230_ (.A(\rbzero.wall_tracer.state[6] ),
    .Y(_04927_));
 sky130_fd_sc_hd__buf_4 _12231_ (.A(_04927_),
    .X(_04928_));
 sky130_fd_sc_hd__buf_4 _12232_ (.A(_04928_),
    .X(_04929_));
 sky130_fd_sc_hd__nor2_1 _12233_ (.A(_04929_),
    .B(_03730_),
    .Y(_00010_));
 sky130_fd_sc_hd__and3_1 _12234_ (.A(o_vsync),
    .B(\rbzero.wall_tracer.state[4] ),
    .C(_03292_),
    .X(_04930_));
 sky130_fd_sc_hd__clkbuf_4 _12235_ (.A(_04930_),
    .X(_04931_));
 sky130_fd_sc_hd__buf_4 _12236_ (.A(_04931_),
    .X(_00008_));
 sky130_fd_sc_hd__inv_2 _12237_ (.A(\rbzero.wall_tracer.state[3] ),
    .Y(_04932_));
 sky130_fd_sc_hd__clkbuf_8 _12238_ (.A(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__nor2_1 _12239_ (.A(_04933_),
    .B(_03730_),
    .Y(_00007_));
 sky130_fd_sc_hd__mux2_1 _12240_ (.A0(\rbzero.debug_overlay.playerY[0] ),
    .A1(_03743_),
    .S(_03798_),
    .X(_04934_));
 sky130_fd_sc_hd__buf_2 _12241_ (.A(\rbzero.wall_tracer.state[6] ),
    .X(_04935_));
 sky130_fd_sc_hd__buf_4 _12242_ (.A(_04935_),
    .X(_04936_));
 sky130_fd_sc_hd__buf_4 _12243_ (.A(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__buf_4 _12244_ (.A(_04937_),
    .X(_04938_));
 sky130_fd_sc_hd__buf_6 _12245_ (.A(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__buf_6 _12246_ (.A(_03731_),
    .X(_04940_));
 sky130_fd_sc_hd__inv_2 _12247_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .Y(_04941_));
 sky130_fd_sc_hd__inv_2 _12248_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .Y(_04942_));
 sky130_fd_sc_hd__o22a_1 _12249_ (.A1(\rbzero.wall_tracer.trackDistX[3] ),
    .A2(_04941_),
    .B1(\rbzero.wall_tracer.trackDistX[2] ),
    .B2(_04942_),
    .X(_04943_));
 sky130_fd_sc_hd__inv_2 _12250_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .Y(_04944_));
 sky130_fd_sc_hd__inv_2 _12251_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .Y(_04945_));
 sky130_fd_sc_hd__o22a_1 _12252_ (.A1(\rbzero.wall_tracer.trackDistX[1] ),
    .A2(_04944_),
    .B1(_04945_),
    .B2(\rbzero.wall_tracer.trackDistX[0] ),
    .X(_04946_));
 sky130_fd_sc_hd__inv_2 _12253_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .Y(_04947_));
 sky130_fd_sc_hd__inv_2 _12254_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .Y(_04948_));
 sky130_fd_sc_hd__a22o_1 _12255_ (.A1(_04947_),
    .A2(\rbzero.wall_tracer.trackDistY[-3] ),
    .B1(\rbzero.wall_tracer.trackDistY[-4] ),
    .B2(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__inv_2 _12256_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .Y(_04950_));
 sky130_fd_sc_hd__o22a_1 _12257_ (.A1(_04950_),
    .A2(\rbzero.wall_tracer.trackDistY[-2] ),
    .B1(_04947_),
    .B2(\rbzero.wall_tracer.trackDistY[-3] ),
    .X(_04951_));
 sky130_fd_sc_hd__nand2_1 _12258_ (.A(_04949_),
    .B(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__inv_2 _12259_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .Y(_04953_));
 sky130_fd_sc_hd__inv_2 _12260_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .Y(_04954_));
 sky130_fd_sc_hd__o22a_1 _12261_ (.A1(\rbzero.wall_tracer.trackDistX[-1] ),
    .A2(_04953_),
    .B1(\rbzero.wall_tracer.trackDistX[-2] ),
    .B2(_04954_),
    .X(_04955_));
 sky130_fd_sc_hd__and2_1 _12262_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(_04953_),
    .X(_04956_));
 sky130_fd_sc_hd__and2_1 _12263_ (.A(_04945_),
    .B(\rbzero.wall_tracer.trackDistX[0] ),
    .X(_04957_));
 sky130_fd_sc_hd__a211o_1 _12264_ (.A1(_04952_),
    .A2(_04955_),
    .B1(_04956_),
    .C1(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__a22o_1 _12265_ (.A1(\rbzero.wall_tracer.trackDistX[2] ),
    .A2(_04942_),
    .B1(\rbzero.wall_tracer.trackDistX[1] ),
    .B2(_04944_),
    .X(_04959_));
 sky130_fd_sc_hd__a21o_1 _12266_ (.A1(_04946_),
    .A2(_04958_),
    .B1(_04959_),
    .X(_04960_));
 sky130_fd_sc_hd__a22o_1 _12267_ (.A1(\rbzero.wall_tracer.trackDistX[3] ),
    .A2(_04941_),
    .B1(_04943_),
    .B2(_04960_),
    .X(_04961_));
 sky130_fd_sc_hd__inv_2 _12268_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .Y(_04962_));
 sky130_fd_sc_hd__inv_2 _12269_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .Y(_04963_));
 sky130_fd_sc_hd__a22o_1 _12270_ (.A1(_04962_),
    .A2(\rbzero.wall_tracer.trackDistY[-7] ),
    .B1(\rbzero.wall_tracer.trackDistY[-8] ),
    .B2(_04963_),
    .X(_04964_));
 sky130_fd_sc_hd__inv_2 _12271_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .Y(_04965_));
 sky130_fd_sc_hd__inv_2 _12272_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .Y(_04966_));
 sky130_fd_sc_hd__or2_1 _12273_ (.A(_04966_),
    .B(\rbzero.wall_tracer.trackDistY[-10] ),
    .X(_04967_));
 sky130_fd_sc_hd__inv_2 _12274_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .Y(_04968_));
 sky130_fd_sc_hd__inv_2 _12275_ (.A(\rbzero.wall_tracer.trackDistX[-12] ),
    .Y(_04969_));
 sky130_fd_sc_hd__o22a_1 _12276_ (.A1(_04968_),
    .A2(\rbzero.wall_tracer.trackDistY[-11] ),
    .B1(\rbzero.wall_tracer.trackDistY[-12] ),
    .B2(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__a21o_1 _12277_ (.A1(_04968_),
    .A2(\rbzero.wall_tracer.trackDistY[-11] ),
    .B1(_04970_),
    .X(_04971_));
 sky130_fd_sc_hd__a22o_1 _12278_ (.A1(_04965_),
    .A2(\rbzero.wall_tracer.trackDistY[-9] ),
    .B1(_04966_),
    .B2(\rbzero.wall_tracer.trackDistY[-10] ),
    .X(_04972_));
 sky130_fd_sc_hd__a21o_1 _12279_ (.A1(_04967_),
    .A2(_04971_),
    .B1(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__o221a_1 _12280_ (.A1(\rbzero.wall_tracer.trackDistY[-8] ),
    .A2(_04963_),
    .B1(_04965_),
    .B2(\rbzero.wall_tracer.trackDistY[-9] ),
    .C1(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__nor2_1 _12281_ (.A(_04964_),
    .B(_04974_),
    .Y(_04975_));
 sky130_fd_sc_hd__nor2_1 _12282_ (.A(_04962_),
    .B(\rbzero.wall_tracer.trackDistY[-7] ),
    .Y(_04976_));
 sky130_fd_sc_hd__inv_2 _12283_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .Y(_04977_));
 sky130_fd_sc_hd__nor2_1 _12284_ (.A(_04977_),
    .B(\rbzero.wall_tracer.trackDistY[-6] ),
    .Y(_04978_));
 sky130_fd_sc_hd__inv_2 _12285_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .Y(_04979_));
 sky130_fd_sc_hd__a22o_1 _12286_ (.A1(_04979_),
    .A2(\rbzero.wall_tracer.trackDistY[-5] ),
    .B1(_04977_),
    .B2(\rbzero.wall_tracer.trackDistY[-6] ),
    .X(_04980_));
 sky130_fd_sc_hd__inv_2 _12287_ (.A(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__o31a_1 _12288_ (.A1(_04975_),
    .A2(_04976_),
    .A3(_04978_),
    .B1(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__nand2_1 _12289_ (.A(_04951_),
    .B(_04955_),
    .Y(_04983_));
 sky130_fd_sc_hd__or4_1 _12290_ (.A(_04956_),
    .B(_04957_),
    .C(_04949_),
    .D(_04983_),
    .X(_04984_));
 sky130_fd_sc_hd__inv_2 _12291_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .Y(_04985_));
 sky130_fd_sc_hd__o221a_1 _12292_ (.A1(_04985_),
    .A2(\rbzero.wall_tracer.trackDistY[3] ),
    .B1(\rbzero.wall_tracer.trackDistY[-4] ),
    .B2(_04948_),
    .C1(_04943_),
    .X(_04986_));
 sky130_fd_sc_hd__nand3b_1 _12293_ (.A_N(_04959_),
    .B(_04946_),
    .C(_04986_),
    .Y(_04987_));
 sky130_fd_sc_hd__or2_1 _12294_ (.A(_04984_),
    .B(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__nor2_1 _12295_ (.A(_04979_),
    .B(\rbzero.wall_tracer.trackDistY[-5] ),
    .Y(_04989_));
 sky130_fd_sc_hd__or3_1 _12296_ (.A(_04982_),
    .B(_04988_),
    .C(_04989_),
    .X(_04990_));
 sky130_fd_sc_hd__inv_2 _12297_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .Y(_04991_));
 sky130_fd_sc_hd__inv_2 _12298_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .Y(_04992_));
 sky130_fd_sc_hd__o22a_1 _12299_ (.A1(\rbzero.wall_tracer.trackDistX[9] ),
    .A2(_04991_),
    .B1(_04992_),
    .B2(\rbzero.wall_tracer.trackDistX[8] ),
    .X(_04993_));
 sky130_fd_sc_hd__inv_2 _12300_ (.A(\rbzero.wall_tracer.trackDistY[11] ),
    .Y(_04994_));
 sky130_fd_sc_hd__inv_2 _12301_ (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .Y(_04995_));
 sky130_fd_sc_hd__o22a_1 _12302_ (.A1(_04994_),
    .A2(\rbzero.wall_tracer.trackDistX[11] ),
    .B1(\rbzero.wall_tracer.trackDistX[10] ),
    .B2(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__nand2_1 _12303_ (.A(_04993_),
    .B(_04996_),
    .Y(_04997_));
 sky130_fd_sc_hd__a22o_1 _12304_ (.A1(\rbzero.wall_tracer.trackDistX[10] ),
    .A2(_04995_),
    .B1(\rbzero.wall_tracer.trackDistX[9] ),
    .B2(_04991_),
    .X(_04998_));
 sky130_fd_sc_hd__inv_2 _12305_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .Y(_04999_));
 sky130_fd_sc_hd__a22o_1 _12306_ (.A1(_04992_),
    .A2(\rbzero.wall_tracer.trackDistX[8] ),
    .B1(\rbzero.wall_tracer.trackDistX[7] ),
    .B2(_04999_),
    .X(_05000_));
 sky130_fd_sc_hd__inv_2 _12307_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .Y(_05001_));
 sky130_fd_sc_hd__inv_2 _12308_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .Y(_05002_));
 sky130_fd_sc_hd__o22a_1 _12309_ (.A1(\rbzero.wall_tracer.trackDistX[5] ),
    .A2(_05002_),
    .B1(_05001_),
    .B2(\rbzero.wall_tracer.trackDistX[4] ),
    .X(_05003_));
 sky130_fd_sc_hd__inv_2 _12310_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .Y(_05004_));
 sky130_fd_sc_hd__o22a_1 _12311_ (.A1(\rbzero.wall_tracer.trackDistX[7] ),
    .A2(_04999_),
    .B1(\rbzero.wall_tracer.trackDistX[6] ),
    .B2(_05004_),
    .X(_05005_));
 sky130_fd_sc_hd__nand2_1 _12312_ (.A(_05003_),
    .B(_05005_),
    .Y(_05006_));
 sky130_fd_sc_hd__a22o_1 _12313_ (.A1(\rbzero.wall_tracer.trackDistX[6] ),
    .A2(_05004_),
    .B1(\rbzero.wall_tracer.trackDistX[5] ),
    .B2(_05002_),
    .X(_05007_));
 sky130_fd_sc_hd__and2_1 _12314_ (.A(_04994_),
    .B(\rbzero.wall_tracer.trackDistX[11] ),
    .X(_05008_));
 sky130_fd_sc_hd__a2111o_1 _12315_ (.A1(_05001_),
    .A2(\rbzero.wall_tracer.trackDistX[4] ),
    .B1(_05006_),
    .C1(_05007_),
    .D1(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__or4_1 _12316_ (.A(_04997_),
    .B(_04998_),
    .C(_05000_),
    .D(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__a21oi_1 _12317_ (.A1(_04961_),
    .A2(_04990_),
    .B1(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__o21a_1 _12318_ (.A1(_05003_),
    .A2(_05007_),
    .B1(_05005_),
    .X(_05012_));
 sky130_fd_sc_hd__o21a_1 _12319_ (.A1(_05000_),
    .A2(_05012_),
    .B1(_04993_),
    .X(_05013_));
 sky130_fd_sc_hd__o21a_1 _12320_ (.A1(_04998_),
    .A2(_05013_),
    .B1(_04996_),
    .X(_05014_));
 sky130_fd_sc_hd__nor2_1 _12321_ (.A(_05008_),
    .B(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__inv_2 _12322_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .Y(_05016_));
 sky130_fd_sc_hd__a211o_1 _12323_ (.A1(_05016_),
    .A2(\rbzero.wall_tracer.trackDistX[-8] ),
    .B1(_04976_),
    .C1(_04978_),
    .X(_05017_));
 sky130_fd_sc_hd__inv_2 _12324_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .Y(_05018_));
 sky130_fd_sc_hd__o21ai_1 _12325_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(_05018_),
    .B1(_04970_),
    .Y(_05019_));
 sky130_fd_sc_hd__inv_2 _12326_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .Y(_05020_));
 sky130_fd_sc_hd__a22o_1 _12327_ (.A1(\rbzero.wall_tracer.trackDistX[-9] ),
    .A2(_05020_),
    .B1(\rbzero.wall_tracer.trackDistY[-12] ),
    .B2(_04969_),
    .X(_05021_));
 sky130_fd_sc_hd__or4b_1 _12328_ (.A(_05019_),
    .B(_04989_),
    .C(_05021_),
    .D_N(_04967_),
    .X(_05022_));
 sky130_fd_sc_hd__or4_1 _12329_ (.A(_04980_),
    .B(_04964_),
    .C(_04972_),
    .D(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__or4_1 _12330_ (.A(_05010_),
    .B(_04988_),
    .C(_05017_),
    .D(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__o21ai_4 _12331_ (.A1(_05011_),
    .A2(_05015_),
    .B1(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__and2_2 _12332_ (.A(_03801_),
    .B(_03779_),
    .X(_05026_));
 sky130_fd_sc_hd__o21a_2 _12333_ (.A1(_04940_),
    .A2(_05025_),
    .B1(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__o21ai_4 _12334_ (.A1(_03798_),
    .A2(_04939_),
    .B1(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__mux2_1 _12335_ (.A0(_04934_),
    .A1(\rbzero.map_rom.d6 ),
    .S(_05028_),
    .X(_05029_));
 sky130_fd_sc_hd__clkbuf_1 _12336_ (.A(_05029_),
    .X(_00401_));
 sky130_fd_sc_hd__xnor2_2 _12337_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_05030_));
 sky130_fd_sc_hd__nand2_1 _12338_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_05031_));
 sky130_fd_sc_hd__or2_1 _12339_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_05032_));
 sky130_fd_sc_hd__nand2_1 _12340_ (.A(_05031_),
    .B(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__nor2_1 _12341_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_05034_));
 sky130_fd_sc_hd__and2_1 _12342_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_05035_));
 sky130_fd_sc_hd__nor2_1 _12343_ (.A(_05034_),
    .B(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__or3b_1 _12344_ (.A(_05030_),
    .B(_05033_),
    .C_N(_05036_),
    .X(_05037_));
 sky130_fd_sc_hd__or2_1 _12345_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_05038_));
 sky130_fd_sc_hd__xor2_2 _12346_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_05039_));
 sky130_fd_sc_hd__and2_1 _12347_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_05040_));
 sky130_fd_sc_hd__a31o_1 _12348_ (.A1(\rbzero.debug_overlay.facingY[-9] ),
    .A2(\rbzero.wall_tracer.rayAddendY[-1] ),
    .A3(_05039_),
    .B1(_05040_),
    .X(_05041_));
 sky130_fd_sc_hd__and2_1 _12349_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_05042_));
 sky130_fd_sc_hd__a221o_1 _12350_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[2] ),
    .B1(_05038_),
    .B2(_05041_),
    .C1(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__or2_1 _12351_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .X(_05044_));
 sky130_fd_sc_hd__nand2_1 _12352_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_05045_));
 sky130_fd_sc_hd__or2_1 _12353_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_05046_));
 sky130_fd_sc_hd__and2_1 _12354_ (.A(_05045_),
    .B(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__and4b_1 _12355_ (.A_N(_05037_),
    .B(_05043_),
    .C(_05044_),
    .D(_05047_),
    .X(_05048_));
 sky130_fd_sc_hd__nand2_1 _12356_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_05049_));
 sky130_fd_sc_hd__a2111oi_1 _12357_ (.A1(_05045_),
    .A2(_05049_),
    .B1(_05034_),
    .C1(_05033_),
    .D1(_05030_),
    .Y(_05050_));
 sky130_fd_sc_hd__o211a_1 _12358_ (.A1(\rbzero.debug_overlay.facingY[-2] ),
    .A2(\rbzero.wall_tracer.rayAddendY[6] ),
    .B1(\rbzero.wall_tracer.rayAddendY[5] ),
    .C1(\rbzero.debug_overlay.facingY[-3] ),
    .X(_05051_));
 sky130_fd_sc_hd__a211o_1 _12359_ (.A1(\rbzero.debug_overlay.facingY[-2] ),
    .A2(\rbzero.wall_tracer.rayAddendY[6] ),
    .B1(_05050_),
    .C1(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__nand2_1 _12360_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .Y(_05053_));
 sky130_fd_sc_hd__or2_1 _12361_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_05054_));
 sky130_fd_sc_hd__and2_1 _12362_ (.A(_05053_),
    .B(_05054_),
    .X(_05055_));
 sky130_fd_sc_hd__o21ai_2 _12363_ (.A1(_05048_),
    .A2(_05052_),
    .B1(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__and2_1 _12364_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .X(_05057_));
 sky130_fd_sc_hd__a21oi_1 _12365_ (.A1(\rbzero.debug_overlay.facingY[-1] ),
    .A2(\rbzero.wall_tracer.rayAddendY[7] ),
    .B1(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__xor2_1 _12366_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .X(_05059_));
 sky130_fd_sc_hd__inv_2 _12367_ (.A(_05059_),
    .Y(_05060_));
 sky130_fd_sc_hd__nand2_1 _12368_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_05061_));
 sky130_fd_sc_hd__or2_1 _12369_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .X(_05062_));
 sky130_fd_sc_hd__nand2_1 _12370_ (.A(_05061_),
    .B(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__nor2_1 _12371_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .Y(_05064_));
 sky130_fd_sc_hd__a2111o_1 _12372_ (.A1(_05056_),
    .A2(_05058_),
    .B1(_05060_),
    .C1(_05063_),
    .D1(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__o21ai_1 _12373_ (.A1(\rbzero.wall_tracer.rayAddendY[10] ),
    .A2(\rbzero.wall_tracer.rayAddendY[9] ),
    .B1(\rbzero.debug_overlay.facingY[10] ),
    .Y(_05066_));
 sky130_fd_sc_hd__nand2_1 _12374_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[11] ),
    .Y(_05067_));
 sky130_fd_sc_hd__or2_1 _12375_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[11] ),
    .X(_05068_));
 sky130_fd_sc_hd__buf_2 _12376_ (.A(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__nand2_1 _12377_ (.A(_05067_),
    .B(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__and3_1 _12378_ (.A(_05065_),
    .B(_05066_),
    .C(_05070_),
    .X(_05071_));
 sky130_fd_sc_hd__a21o_1 _12379_ (.A1(_05065_),
    .A2(_05066_),
    .B1(_05070_),
    .X(_05072_));
 sky130_fd_sc_hd__and2b_1 _12380_ (.A_N(_05071_),
    .B(_05072_),
    .X(_05073_));
 sky130_fd_sc_hd__nand3_1 _12381_ (.A(_05044_),
    .B(_05043_),
    .C(_05047_),
    .Y(_05074_));
 sky130_fd_sc_hd__a311o_2 _12382_ (.A1(_05045_),
    .A2(_05074_),
    .A3(_05049_),
    .B1(_05034_),
    .C1(_05033_),
    .X(_05075_));
 sky130_fd_sc_hd__a21o_1 _12383_ (.A1(_05031_),
    .A2(_05075_),
    .B1(_05030_),
    .X(_05076_));
 sky130_fd_sc_hd__nand3_1 _12384_ (.A(_05030_),
    .B(_05031_),
    .C(_05075_),
    .Y(_05077_));
 sky130_fd_sc_hd__and2_1 _12385_ (.A(_05076_),
    .B(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__a21oi_1 _12386_ (.A1(_05056_),
    .A2(_05058_),
    .B1(_05064_),
    .Y(_05079_));
 sky130_fd_sc_hd__xnor2_2 _12387_ (.A(_05063_),
    .B(_05079_),
    .Y(_05080_));
 sky130_fd_sc_hd__inv_2 _12388_ (.A(_05034_),
    .Y(_05081_));
 sky130_fd_sc_hd__a32o_1 _12389_ (.A1(_05044_),
    .A2(_05043_),
    .A3(_05047_),
    .B1(\rbzero.wall_tracer.rayAddendY[3] ),
    .B2(\rbzero.debug_overlay.facingY[-5] ),
    .X(_05082_));
 sky130_fd_sc_hd__a221o_1 _12390_ (.A1(_05031_),
    .A2(_05032_),
    .B1(_05081_),
    .B2(_05082_),
    .C1(_05035_),
    .X(_05083_));
 sky130_fd_sc_hd__and2_1 _12391_ (.A(_05075_),
    .B(_05083_),
    .X(_05084_));
 sky130_fd_sc_hd__xor2_2 _12392_ (.A(_05036_),
    .B(_05082_),
    .X(_05085_));
 sky130_fd_sc_hd__nand2_1 _12393_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_05086_));
 sky130_fd_sc_hd__nand2_1 _12394_ (.A(_05044_),
    .B(_05086_),
    .Y(_05087_));
 sky130_fd_sc_hd__a21o_1 _12395_ (.A1(_05038_),
    .A2(_05041_),
    .B1(_05042_),
    .X(_05088_));
 sky130_fd_sc_hd__xnor2_2 _12396_ (.A(_05087_),
    .B(_05088_),
    .Y(_05089_));
 sky130_fd_sc_hd__a21o_1 _12397_ (.A1(_05044_),
    .A2(_05043_),
    .B1(_05047_),
    .X(_05090_));
 sky130_fd_sc_hd__and2_1 _12398_ (.A(_05074_),
    .B(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__or2b_1 _12399_ (.A(_05042_),
    .B_N(_05038_),
    .X(_05092_));
 sky130_fd_sc_hd__xnor2_2 _12400_ (.A(_05092_),
    .B(_05041_),
    .Y(_05093_));
 sky130_fd_sc_hd__nand2_1 _12401_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_05094_));
 sky130_fd_sc_hd__xnor2_2 _12402_ (.A(_05094_),
    .B(_05039_),
    .Y(_05095_));
 sky130_fd_sc_hd__xor2_2 _12403_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_05096_));
 sky130_fd_sc_hd__or4_1 _12404_ (.A(\rbzero.wall_tracer.rayAddendY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .C(_05095_),
    .D(_05096_),
    .X(_05097_));
 sky130_fd_sc_hd__or4_1 _12405_ (.A(\rbzero.wall_tracer.rayAddendY[-4] ),
    .B(_05091_),
    .C(_05093_),
    .D(_05097_),
    .X(_05098_));
 sky130_fd_sc_hd__or3_1 _12406_ (.A(_05055_),
    .B(_05048_),
    .C(_05052_),
    .X(_05099_));
 sky130_fd_sc_hd__and2_1 _12407_ (.A(_05056_),
    .B(_05099_),
    .X(_05100_));
 sky130_fd_sc_hd__or4_1 _12408_ (.A(_05085_),
    .B(_05089_),
    .C(_05098_),
    .D(_05100_),
    .X(_05101_));
 sky130_fd_sc_hd__or4_1 _12409_ (.A(_05078_),
    .B(_05080_),
    .C(_05084_),
    .D(_05101_),
    .X(_05102_));
 sky130_fd_sc_hd__a211o_1 _12410_ (.A1(_05056_),
    .A2(_05058_),
    .B1(_05063_),
    .C1(_05064_),
    .X(_05103_));
 sky130_fd_sc_hd__nand3_1 _12411_ (.A(_05059_),
    .B(_05061_),
    .C(_05103_),
    .Y(_05104_));
 sky130_fd_sc_hd__a21o_1 _12412_ (.A1(_05061_),
    .A2(_05103_),
    .B1(_05059_),
    .X(_05105_));
 sky130_fd_sc_hd__nand2_1 _12413_ (.A(_05104_),
    .B(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__nor2_1 _12414_ (.A(_05064_),
    .B(_05057_),
    .Y(_05107_));
 sky130_fd_sc_hd__a21oi_1 _12415_ (.A1(_05053_),
    .A2(_05056_),
    .B1(_05107_),
    .Y(_05108_));
 sky130_fd_sc_hd__and3_1 _12416_ (.A(_05053_),
    .B(_05056_),
    .C(_05107_),
    .X(_05109_));
 sky130_fd_sc_hd__nor2_1 _12417_ (.A(_05108_),
    .B(_05109_),
    .Y(_05110_));
 sky130_fd_sc_hd__or3b_1 _12418_ (.A(_05102_),
    .B(_05106_),
    .C_N(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__a21bo_2 _12419_ (.A1(_05065_),
    .A2(_05066_),
    .B1_N(_05067_),
    .X(_05112_));
 sky130_fd_sc_hd__a2bb2o_4 _12420_ (.A1_N(_05073_),
    .A2_N(_05111_),
    .B1(_05112_),
    .B2(_05069_),
    .X(_05113_));
 sky130_fd_sc_hd__buf_4 _12421_ (.A(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__and2_1 _12422_ (.A(\rbzero.map_rom.c6 ),
    .B(_05114_),
    .X(_05115_));
 sky130_fd_sc_hd__nor2_1 _12423_ (.A(\rbzero.map_rom.c6 ),
    .B(_05114_),
    .Y(_05116_));
 sky130_fd_sc_hd__nor2_1 _12424_ (.A(_05115_),
    .B(_05116_),
    .Y(_05117_));
 sky130_fd_sc_hd__xnor2_1 _12425_ (.A(_03743_),
    .B(_05117_),
    .Y(_05118_));
 sky130_fd_sc_hd__mux2_1 _12426_ (.A0(\rbzero.debug_overlay.playerY[1] ),
    .A1(_05118_),
    .S(_03798_),
    .X(_05119_));
 sky130_fd_sc_hd__mux2_1 _12427_ (.A0(_05119_),
    .A1(\rbzero.map_rom.c6 ),
    .S(_05028_),
    .X(_05120_));
 sky130_fd_sc_hd__clkbuf_1 _12428_ (.A(_05120_),
    .X(_00402_));
 sky130_fd_sc_hd__buf_6 _12429_ (.A(_03797_),
    .X(_05121_));
 sky130_fd_sc_hd__nand2_1 _12430_ (.A(_03733_),
    .B(_05114_),
    .Y(_05122_));
 sky130_fd_sc_hd__or2_1 _12431_ (.A(_03733_),
    .B(_05114_),
    .X(_05123_));
 sky130_fd_sc_hd__and2_1 _12432_ (.A(_05122_),
    .B(_05123_),
    .X(_05124_));
 sky130_fd_sc_hd__a21o_1 _12433_ (.A1(\rbzero.map_rom.d6 ),
    .A2(_05117_),
    .B1(_05115_),
    .X(_05125_));
 sky130_fd_sc_hd__or2_1 _12434_ (.A(_05124_),
    .B(_05125_),
    .X(_05126_));
 sky130_fd_sc_hd__nand2_1 _12435_ (.A(_05124_),
    .B(_05125_),
    .Y(_05127_));
 sky130_fd_sc_hd__and2_1 _12436_ (.A(\rbzero.debug_overlay.playerY[2] ),
    .B(_04940_),
    .X(_05128_));
 sky130_fd_sc_hd__a31o_1 _12437_ (.A1(_05121_),
    .A2(_05126_),
    .A3(_05127_),
    .B1(_05128_),
    .X(_05129_));
 sky130_fd_sc_hd__mux2_1 _12438_ (.A0(_05129_),
    .A1(_03733_),
    .S(_05028_),
    .X(_05130_));
 sky130_fd_sc_hd__clkbuf_1 _12439_ (.A(_05130_),
    .X(_00403_));
 sky130_fd_sc_hd__nand2_1 _12440_ (.A(\rbzero.map_rom.a6 ),
    .B(_05114_),
    .Y(_05131_));
 sky130_fd_sc_hd__or2_1 _12441_ (.A(\rbzero.map_rom.a6 ),
    .B(_05114_),
    .X(_05132_));
 sky130_fd_sc_hd__nand2_1 _12442_ (.A(_05131_),
    .B(_05132_),
    .Y(_05133_));
 sky130_fd_sc_hd__nand2_1 _12443_ (.A(_05122_),
    .B(_05127_),
    .Y(_05134_));
 sky130_fd_sc_hd__xnor2_1 _12444_ (.A(_05133_),
    .B(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__mux2_1 _12445_ (.A0(\rbzero.debug_overlay.playerY[3] ),
    .A1(_05135_),
    .S(_03798_),
    .X(_05136_));
 sky130_fd_sc_hd__mux2_1 _12446_ (.A0(_05136_),
    .A1(\rbzero.map_rom.a6 ),
    .S(_05028_),
    .X(_05137_));
 sky130_fd_sc_hd__clkbuf_1 _12447_ (.A(_05137_),
    .X(_00404_));
 sky130_fd_sc_hd__xnor2_1 _12448_ (.A(_03732_),
    .B(_05114_),
    .Y(_05138_));
 sky130_fd_sc_hd__o211a_1 _12449_ (.A1(_05127_),
    .A2(_05133_),
    .B1(_05131_),
    .C1(_05122_),
    .X(_05139_));
 sky130_fd_sc_hd__xnor2_1 _12450_ (.A(_05138_),
    .B(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__mux2_1 _12451_ (.A0(\rbzero.debug_overlay.playerY[4] ),
    .A1(_05140_),
    .S(_03798_),
    .X(_05141_));
 sky130_fd_sc_hd__mux2_1 _12452_ (.A0(_05141_),
    .A1(\rbzero.map_rom.i_row[4] ),
    .S(_05028_),
    .X(_05142_));
 sky130_fd_sc_hd__clkbuf_1 _12453_ (.A(_05142_),
    .X(_00405_));
 sky130_fd_sc_hd__nand2_2 _12454_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[11] ),
    .Y(_05143_));
 sky130_fd_sc_hd__or2_1 _12455_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .X(_05144_));
 sky130_fd_sc_hd__and2_1 _12456_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .X(_05145_));
 sky130_fd_sc_hd__a31o_1 _12457_ (.A1(\rbzero.debug_overlay.facingX[-1] ),
    .A2(\rbzero.wall_tracer.rayAddendX[7] ),
    .A3(_05144_),
    .B1(_05145_),
    .X(_05146_));
 sky130_fd_sc_hd__nor2_1 _12458_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_05147_));
 sky130_fd_sc_hd__nor2_1 _12459_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_05148_));
 sky130_fd_sc_hd__nand2_2 _12460_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_05149_));
 sky130_fd_sc_hd__nor2_1 _12461_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_05150_));
 sky130_fd_sc_hd__nand2_1 _12462_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_05151_));
 sky130_fd_sc_hd__nand2_1 _12463_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_05152_));
 sky130_fd_sc_hd__o211a_1 _12464_ (.A1(_05149_),
    .A2(_05150_),
    .B1(_05151_),
    .C1(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__nand2_1 _12465_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_05154_));
 sky130_fd_sc_hd__o31a_2 _12466_ (.A1(_05147_),
    .A2(_05148_),
    .A3(_05153_),
    .B1(_05154_),
    .X(_05155_));
 sky130_fd_sc_hd__nand2_1 _12467_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_05156_));
 sky130_fd_sc_hd__or2_1 _12468_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_05157_));
 sky130_fd_sc_hd__nand2_2 _12469_ (.A(_05156_),
    .B(_05157_),
    .Y(_05158_));
 sky130_fd_sc_hd__or2_1 _12470_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .X(_05159_));
 sky130_fd_sc_hd__nand2_1 _12471_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .Y(_05160_));
 sky130_fd_sc_hd__and2_1 _12472_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_05161_));
 sky130_fd_sc_hd__nor2_1 _12473_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_05162_));
 sky130_fd_sc_hd__nor2_2 _12474_ (.A(_05161_),
    .B(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__and3_1 _12475_ (.A(_05159_),
    .B(_05160_),
    .C(_05163_),
    .X(_05164_));
 sky130_fd_sc_hd__nor2_1 _12476_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .Y(_05165_));
 sky130_fd_sc_hd__nand2_1 _12477_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .Y(_05166_));
 sky130_fd_sc_hd__and2b_1 _12478_ (.A_N(_05165_),
    .B(_05166_),
    .X(_05167_));
 sky130_fd_sc_hd__and4bb_1 _12479_ (.A_N(_05155_),
    .B_N(_05158_),
    .C(_05164_),
    .D(_05167_),
    .X(_05168_));
 sky130_fd_sc_hd__a21oi_1 _12480_ (.A1(_05156_),
    .A2(_05166_),
    .B1(_05165_),
    .Y(_05169_));
 sky130_fd_sc_hd__and2_1 _12481_ (.A(_05159_),
    .B(_05161_),
    .X(_05170_));
 sky130_fd_sc_hd__a221o_1 _12482_ (.A1(\rbzero.debug_overlay.facingX[-2] ),
    .A2(\rbzero.wall_tracer.rayAddendX[6] ),
    .B1(_05164_),
    .B2(_05169_),
    .C1(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__or2b_1 _12483_ (.A(_05145_),
    .B_N(_05144_),
    .X(_05172_));
 sky130_fd_sc_hd__inv_2 _12484_ (.A(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__nand2_1 _12485_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .Y(_05174_));
 sky130_fd_sc_hd__or2_1 _12486_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_05175_));
 sky130_fd_sc_hd__and2_1 _12487_ (.A(_05174_),
    .B(_05175_),
    .X(_05176_));
 sky130_fd_sc_hd__o211a_1 _12488_ (.A1(_05168_),
    .A2(_05171_),
    .B1(_05173_),
    .C1(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__or2_1 _12489_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_05178_));
 sky130_fd_sc_hd__nand2_1 _12490_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_05179_));
 sky130_fd_sc_hd__nand2_2 _12491_ (.A(_05178_),
    .B(_05179_),
    .Y(_05180_));
 sky130_fd_sc_hd__o21bai_1 _12492_ (.A1(_05146_),
    .A2(_05177_),
    .B1_N(_05180_),
    .Y(_05181_));
 sky130_fd_sc_hd__xnor2_2 _12493_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_05182_));
 sky130_fd_sc_hd__or2_1 _12494_ (.A(\rbzero.wall_tracer.rayAddendX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_05183_));
 sky130_fd_sc_hd__a2bb2o_4 _12495_ (.A1_N(_05181_),
    .A2_N(_05182_),
    .B1(\rbzero.debug_overlay.facingX[10] ),
    .B2(_05183_),
    .X(_05184_));
 sky130_fd_sc_hd__nor2_2 _12496_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[11] ),
    .Y(_05185_));
 sky130_fd_sc_hd__a21oi_4 _12497_ (.A1(_05143_),
    .A2(_05184_),
    .B1(_05185_),
    .Y(_05186_));
 sky130_fd_sc_hd__nand2_1 _12498_ (.A(_03790_),
    .B(_05186_),
    .Y(_05187_));
 sky130_fd_sc_hd__nand3_2 _12499_ (.A(_03816_),
    .B(_05069_),
    .C(_05112_),
    .Y(_05188_));
 sky130_fd_sc_hd__inv_2 _12500_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .Y(_05189_));
 sky130_fd_sc_hd__buf_2 _12501_ (.A(_05189_),
    .X(_05190_));
 sky130_fd_sc_hd__nand2_1 _12502_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__a21o_1 _12503_ (.A1(_05188_),
    .A2(_05191_),
    .B1(_03790_),
    .X(_05192_));
 sky130_fd_sc_hd__nand2_1 _12504_ (.A(_05187_),
    .B(_05192_),
    .Y(_05193_));
 sky130_fd_sc_hd__or2_1 _12505_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[11] ),
    .X(_05194_));
 sky130_fd_sc_hd__nand2_1 _12506_ (.A(_05143_),
    .B(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__xor2_2 _12507_ (.A(_05184_),
    .B(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__a21o_1 _12508_ (.A1(\rbzero.wall_tracer.visualWallDist[3] ),
    .A2(_05190_),
    .B1(_03789_),
    .X(_05197_));
 sky130_fd_sc_hd__and3b_1 _12509_ (.A_N(_05071_),
    .B(_05072_),
    .C(_03815_),
    .X(_05198_));
 sky130_fd_sc_hd__o2bb2a_2 _12510_ (.A1_N(_03789_),
    .A2_N(_05196_),
    .B1(_05197_),
    .B2(_05198_),
    .X(_05199_));
 sky130_fd_sc_hd__nand2_1 _12511_ (.A(_03816_),
    .B(_05080_),
    .Y(_05200_));
 sky130_fd_sc_hd__a21oi_2 _12512_ (.A1(\rbzero.wall_tracer.visualWallDist[1] ),
    .A2(_05190_),
    .B1(_03789_),
    .Y(_05201_));
 sky130_fd_sc_hd__nor2_2 _12513_ (.A(_05146_),
    .B(_05177_),
    .Y(_05202_));
 sky130_fd_sc_hd__xnor2_4 _12514_ (.A(_05180_),
    .B(_05202_),
    .Y(_05203_));
 sky130_fd_sc_hd__a22oi_4 _12515_ (.A1(_05200_),
    .A2(_05201_),
    .B1(_05203_),
    .B2(_03789_),
    .Y(_05204_));
 sky130_fd_sc_hd__nand2_1 _12516_ (.A(_05159_),
    .B(_05160_),
    .Y(_05205_));
 sky130_fd_sc_hd__inv_2 _12517_ (.A(_05167_),
    .Y(_05206_));
 sky130_fd_sc_hd__inv_2 _12518_ (.A(_05169_),
    .Y(_05207_));
 sky130_fd_sc_hd__o31a_2 _12519_ (.A1(_05155_),
    .A2(_05158_),
    .A3(_05206_),
    .B1(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__o21ba_1 _12520_ (.A1(_05162_),
    .A2(_05208_),
    .B1_N(_05161_),
    .X(_05209_));
 sky130_fd_sc_hd__xnor2_2 _12521_ (.A(_05205_),
    .B(_05209_),
    .Y(_05210_));
 sky130_fd_sc_hd__nand2_1 _12522_ (.A(_03789_),
    .B(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__a21o_1 _12523_ (.A1(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A2(_05190_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_05212_));
 sky130_fd_sc_hd__a31o_1 _12524_ (.A1(_03815_),
    .A2(_05076_),
    .A3(_05077_),
    .B1(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__or2_1 _12525_ (.A(_05168_),
    .B(_05171_),
    .X(_05214_));
 sky130_fd_sc_hd__xnor2_2 _12526_ (.A(_05176_),
    .B(_05214_),
    .Y(_05215_));
 sky130_fd_sc_hd__and3_1 _12527_ (.A(_03815_),
    .B(_05056_),
    .C(_05099_),
    .X(_05216_));
 sky130_fd_sc_hd__a21o_1 _12528_ (.A1(\rbzero.wall_tracer.visualWallDist[-1] ),
    .A2(_05189_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_05217_));
 sky130_fd_sc_hd__o2bb2a_2 _12529_ (.A1_N(_03789_),
    .A2_N(_05215_),
    .B1(_05216_),
    .B2(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__inv_2 _12530_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .Y(_05219_));
 sky130_fd_sc_hd__buf_4 _12531_ (.A(_05219_),
    .X(_05220_));
 sky130_fd_sc_hd__xnor2_4 _12532_ (.A(_05163_),
    .B(_05208_),
    .Y(_05221_));
 sky130_fd_sc_hd__a21o_1 _12533_ (.A1(\rbzero.wall_tracer.visualWallDist[-3] ),
    .A2(_05189_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_05222_));
 sky130_fd_sc_hd__a31o_1 _12534_ (.A1(_03815_),
    .A2(_05075_),
    .A3(_05083_),
    .B1(_05222_),
    .X(_05223_));
 sky130_fd_sc_hd__o21a_1 _12535_ (.A1(_05220_),
    .A2(_05221_),
    .B1(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__o21a_1 _12536_ (.A1(_05155_),
    .A2(_05158_),
    .B1(_05156_),
    .X(_05225_));
 sky130_fd_sc_hd__xnor2_2 _12537_ (.A(_05167_),
    .B(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__or2_1 _12538_ (.A(_05219_),
    .B(_05226_),
    .X(_05227_));
 sky130_fd_sc_hd__a21o_1 _12539_ (.A1(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A2(_05189_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_05228_));
 sky130_fd_sc_hd__a21o_1 _12540_ (.A1(_03815_),
    .A2(_05085_),
    .B1(_05228_),
    .X(_05229_));
 sky130_fd_sc_hd__xnor2_2 _12541_ (.A(_05155_),
    .B(_05158_),
    .Y(_05230_));
 sky130_fd_sc_hd__a21o_1 _12542_ (.A1(\rbzero.wall_tracer.visualWallDist[-5] ),
    .A2(_05189_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_05231_));
 sky130_fd_sc_hd__and3_1 _12543_ (.A(_03815_),
    .B(_05074_),
    .C(_05090_),
    .X(_05232_));
 sky130_fd_sc_hd__o2bb2a_1 _12544_ (.A1_N(\rbzero.wall_tracer.rcp_sel[0] ),
    .A2_N(_05230_),
    .B1(_05231_),
    .B2(_05232_),
    .X(_05233_));
 sky130_fd_sc_hd__nor2_1 _12545_ (.A(_05148_),
    .B(_05153_),
    .Y(_05234_));
 sky130_fd_sc_hd__or2b_1 _12546_ (.A(_05147_),
    .B_N(_05154_),
    .X(_05235_));
 sky130_fd_sc_hd__xnor2_2 _12547_ (.A(_05234_),
    .B(_05235_),
    .Y(_05236_));
 sky130_fd_sc_hd__or2_1 _12548_ (.A(_05219_),
    .B(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__a21o_1 _12549_ (.A1(\rbzero.wall_tracer.visualWallDist[-6] ),
    .A2(_05189_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_05238_));
 sky130_fd_sc_hd__a21o_1 _12550_ (.A1(_03815_),
    .A2(_05089_),
    .B1(_05238_),
    .X(_05239_));
 sky130_fd_sc_hd__o21a_1 _12551_ (.A1(_05149_),
    .A2(_05150_),
    .B1(_05152_),
    .X(_05240_));
 sky130_fd_sc_hd__and2b_1 _12552_ (.A_N(_05148_),
    .B(_05151_),
    .X(_05241_));
 sky130_fd_sc_hd__xnor2_4 _12553_ (.A(_05240_),
    .B(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__or2_1 _12554_ (.A(\rbzero.wall_tracer.visualWallDist[-7] ),
    .B(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05243_));
 sky130_fd_sc_hd__o211a_1 _12555_ (.A1(_05189_),
    .A2(_05093_),
    .B1(_05243_),
    .C1(_05219_),
    .X(_05244_));
 sky130_fd_sc_hd__and2_1 _12556_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_05245_));
 sky130_fd_sc_hd__nor2_1 _12557_ (.A(_05245_),
    .B(_05150_),
    .Y(_05246_));
 sky130_fd_sc_hd__xnor2_2 _12558_ (.A(_05149_),
    .B(_05246_),
    .Y(_05247_));
 sky130_fd_sc_hd__mux2_1 _12559_ (.A0(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A1(_05095_),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05248_));
 sky130_fd_sc_hd__mux2_2 _12560_ (.A0(_05247_),
    .A1(_05248_),
    .S(_05219_),
    .X(_05249_));
 sky130_fd_sc_hd__mux2_1 _12561_ (.A0(\rbzero.wall_tracer.visualWallDist[-10] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-2] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05250_));
 sky130_fd_sc_hd__mux2_2 _12562_ (.A0(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A1(_05250_),
    .S(_05219_),
    .X(_05251_));
 sky130_fd_sc_hd__mux2_1 _12563_ (.A0(\rbzero.wall_tracer.visualWallDist[-12] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-4] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05252_));
 sky130_fd_sc_hd__mux2_4 _12564_ (.A0(\rbzero.wall_tracer.rayAddendX[-4] ),
    .A1(_05252_),
    .S(_05219_),
    .X(_05253_));
 sky130_fd_sc_hd__mux2_1 _12565_ (.A0(\rbzero.wall_tracer.visualWallDist[-11] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-3] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05254_));
 sky130_fd_sc_hd__mux2_2 _12566_ (.A0(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A1(_05254_),
    .S(_05219_),
    .X(_05255_));
 sky130_fd_sc_hd__or3_1 _12567_ (.A(_05251_),
    .B(_05253_),
    .C(_05255_),
    .X(_05256_));
 sky130_fd_sc_hd__or2_1 _12568_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_05257_));
 sky130_fd_sc_hd__and2_1 _12569_ (.A(_05149_),
    .B(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__mux2_1 _12570_ (.A0(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A1(_05096_),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05259_));
 sky130_fd_sc_hd__mux2_2 _12571_ (.A0(_05258_),
    .A1(_05259_),
    .S(_05219_),
    .X(_05260_));
 sky130_fd_sc_hd__or2_1 _12572_ (.A(_05256_),
    .B(_05260_),
    .X(_05261_));
 sky130_fd_sc_hd__a2111o_1 _12573_ (.A1(\rbzero.wall_tracer.rcp_sel[0] ),
    .A2(_05242_),
    .B1(_05244_),
    .C1(_05249_),
    .D1(_05261_),
    .X(_05262_));
 sky130_fd_sc_hd__a21o_1 _12574_ (.A1(_05237_),
    .A2(_05239_),
    .B1(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__a211o_1 _12575_ (.A1(_05227_),
    .A2(_05229_),
    .B1(_05233_),
    .C1(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__a2111o_1 _12576_ (.A1(_05211_),
    .A2(_05213_),
    .B1(_05218_),
    .C1(_05224_),
    .D1(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__a21bo_1 _12577_ (.A1(_05175_),
    .A2(_05214_),
    .B1_N(_05174_),
    .X(_05266_));
 sky130_fd_sc_hd__xnor2_2 _12578_ (.A(_05266_),
    .B(_05172_),
    .Y(_05267_));
 sky130_fd_sc_hd__o21ai_1 _12579_ (.A1(_05108_),
    .A2(_05109_),
    .B1(_03815_),
    .Y(_05268_));
 sky130_fd_sc_hd__a21oi_1 _12580_ (.A1(\rbzero.wall_tracer.visualWallDist[0] ),
    .A2(_05190_),
    .B1(_03789_),
    .Y(_05269_));
 sky130_fd_sc_hd__a2bb2o_1 _12581_ (.A1_N(_05220_),
    .A2_N(_05267_),
    .B1(_05268_),
    .B2(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__nand2b_1 _12582_ (.A_N(_05265_),
    .B(_05270_),
    .Y(_05271_));
 sky130_fd_sc_hd__nand2_1 _12583_ (.A(_05179_),
    .B(_05181_),
    .Y(_05272_));
 sky130_fd_sc_hd__xnor2_2 _12584_ (.A(_05182_),
    .B(_05272_),
    .Y(_05273_));
 sky130_fd_sc_hd__nor2_1 _12585_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_03815_),
    .Y(_05274_));
 sky130_fd_sc_hd__a311o_1 _12586_ (.A1(_03816_),
    .A2(_05104_),
    .A3(_05105_),
    .B1(_05274_),
    .C1(_03789_),
    .X(_05275_));
 sky130_fd_sc_hd__a21bo_2 _12587_ (.A1(_03789_),
    .A2(_05273_),
    .B1_N(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__or4_2 _12588_ (.A(_05199_),
    .B(_05204_),
    .C(_05271_),
    .D(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__and2_1 _12589_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_05190_),
    .X(_05278_));
 sky130_fd_sc_hd__a31o_1 _12590_ (.A1(_03816_),
    .A2(_05069_),
    .A3(_05112_),
    .B1(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__a211oi_4 _12591_ (.A1(_05143_),
    .A2(_05184_),
    .B1(_05185_),
    .C1(_05220_),
    .Y(_05280_));
 sky130_fd_sc_hd__a21o_1 _12592_ (.A1(_05220_),
    .A2(_05279_),
    .B1(_05280_),
    .X(_05281_));
 sky130_fd_sc_hd__and2_1 _12593_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_05190_),
    .X(_05282_));
 sky130_fd_sc_hd__a31o_1 _12594_ (.A1(_03816_),
    .A2(_05069_),
    .A3(_05112_),
    .B1(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__a21o_1 _12595_ (.A1(_05220_),
    .A2(_05283_),
    .B1(_05280_),
    .X(_05284_));
 sky130_fd_sc_hd__nand2_1 _12596_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_05190_),
    .Y(_05285_));
 sky130_fd_sc_hd__a21oi_1 _12597_ (.A1(_05188_),
    .A2(_05285_),
    .B1(_03790_),
    .Y(_05286_));
 sky130_fd_sc_hd__nand2_1 _12598_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_05190_),
    .Y(_05287_));
 sky130_fd_sc_hd__a21o_1 _12599_ (.A1(_05188_),
    .A2(_05287_),
    .B1(_03790_),
    .X(_05288_));
 sky130_fd_sc_hd__or4b_2 _12600_ (.A(_05281_),
    .B(_05284_),
    .C(_05286_),
    .D_N(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__clkinv_2 _12601_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .Y(_05290_));
 sky130_fd_sc_hd__o21a_1 _12602_ (.A1(_05290_),
    .A2(_03816_),
    .B1(_05188_),
    .X(_05291_));
 sky130_fd_sc_hd__o21ai_2 _12603_ (.A1(_03790_),
    .A2(_05291_),
    .B1(_05187_),
    .Y(_05292_));
 sky130_fd_sc_hd__and2_1 _12604_ (.A(\rbzero.wall_tracer.visualWallDist[11] ),
    .B(_05190_),
    .X(_05293_));
 sky130_fd_sc_hd__a31o_1 _12605_ (.A1(_03816_),
    .A2(_05069_),
    .A3(_05112_),
    .B1(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__a21o_1 _12606_ (.A1(_05220_),
    .A2(_05294_),
    .B1(_05280_),
    .X(_05295_));
 sky130_fd_sc_hd__buf_2 _12607_ (.A(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__o31a_1 _12608_ (.A1(_05277_),
    .A2(_05289_),
    .A3(_05292_),
    .B1(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__xnor2_2 _12609_ (.A(_05193_),
    .B(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__o21a_1 _12610_ (.A1(_05277_),
    .A2(_05289_),
    .B1(_05296_),
    .X(_05299_));
 sky130_fd_sc_hd__xnor2_1 _12611_ (.A(_05292_),
    .B(_05299_),
    .Y(_05300_));
 sky130_fd_sc_hd__clkinv_2 _12612_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .Y(_05301_));
 sky130_fd_sc_hd__o21ai_1 _12613_ (.A1(_05301_),
    .A2(_03816_),
    .B1(_05188_),
    .Y(_05302_));
 sky130_fd_sc_hd__a21o_1 _12614_ (.A1(_05220_),
    .A2(_05302_),
    .B1(_05280_),
    .X(_05303_));
 sky130_fd_sc_hd__o211ai_1 _12615_ (.A1(_03790_),
    .A2(_05291_),
    .B1(_05192_),
    .C1(_05187_),
    .Y(_05304_));
 sky130_fd_sc_hd__clkbuf_4 _12616_ (.A(_05296_),
    .X(_05305_));
 sky130_fd_sc_hd__o31a_1 _12617_ (.A1(_05277_),
    .A2(_05289_),
    .A3(_05304_),
    .B1(_05305_),
    .X(_05306_));
 sky130_fd_sc_hd__xnor2_1 _12618_ (.A(_05303_),
    .B(_05306_),
    .Y(_05307_));
 sky130_fd_sc_hd__or4b_1 _12619_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_03816_),
    .C(_03790_),
    .D_N(\rbzero.wall_tracer.visualWallDist[11] ),
    .X(_05308_));
 sky130_fd_sc_hd__or4_1 _12620_ (.A(_05277_),
    .B(_05289_),
    .C(_05304_),
    .D(_05308_),
    .X(_05309_));
 sky130_fd_sc_hd__and4_1 _12621_ (.A(_05298_),
    .B(_05300_),
    .C(_05307_),
    .D(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__a21oi_2 _12622_ (.A1(_05220_),
    .A2(_05283_),
    .B1(_05280_),
    .Y(_05311_));
 sky130_fd_sc_hd__nand2_1 _12623_ (.A(_05288_),
    .B(_05311_),
    .Y(_05312_));
 sky130_fd_sc_hd__o31ai_2 _12624_ (.A1(_05277_),
    .A2(_05312_),
    .A3(_05286_),
    .B1(_05305_),
    .Y(_05313_));
 sky130_fd_sc_hd__xnor2_2 _12625_ (.A(_05281_),
    .B(_05313_),
    .Y(_05314_));
 sky130_fd_sc_hd__nor2_1 _12626_ (.A(_05280_),
    .B(_05286_),
    .Y(_05315_));
 sky130_fd_sc_hd__o41a_2 _12627_ (.A1(_05199_),
    .A2(_05204_),
    .A3(_05271_),
    .A4(_05276_),
    .B1(_05296_),
    .X(_05316_));
 sky130_fd_sc_hd__a21o_1 _12628_ (.A1(_05305_),
    .A2(_05312_),
    .B1(_05316_),
    .X(_05317_));
 sky130_fd_sc_hd__xor2_1 _12629_ (.A(_05315_),
    .B(_05317_),
    .X(_05318_));
 sky130_fd_sc_hd__nand2_1 _12630_ (.A(_05187_),
    .B(_05288_),
    .Y(_05319_));
 sky130_fd_sc_hd__a21o_1 _12631_ (.A1(_05305_),
    .A2(_05284_),
    .B1(_05316_),
    .X(_05320_));
 sky130_fd_sc_hd__xnor2_2 _12632_ (.A(_05319_),
    .B(_05320_),
    .Y(_05321_));
 sky130_fd_sc_hd__and3b_1 _12633_ (.A_N(_05314_),
    .B(_05318_),
    .C(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__xnor2_2 _12634_ (.A(_05311_),
    .B(_05316_),
    .Y(_05323_));
 sky130_fd_sc_hd__o31a_1 _12635_ (.A1(_05204_),
    .A2(_05271_),
    .A3(_05276_),
    .B1(_05296_),
    .X(_05324_));
 sky130_fd_sc_hd__xor2_4 _12636_ (.A(_05199_),
    .B(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__o21ai_1 _12637_ (.A1(_05204_),
    .A2(_05271_),
    .B1(_05305_),
    .Y(_05326_));
 sky130_fd_sc_hd__xnor2_2 _12638_ (.A(_05276_),
    .B(_05326_),
    .Y(_05327_));
 sky130_fd_sc_hd__or2_1 _12639_ (.A(_05325_),
    .B(_05327_),
    .X(_05328_));
 sky130_fd_sc_hd__nor2_1 _12640_ (.A(_05323_),
    .B(_05328_),
    .Y(_05329_));
 sky130_fd_sc_hd__a22o_1 _12641_ (.A1(_05200_),
    .A2(_05201_),
    .B1(_05203_),
    .B2(_03790_),
    .X(_05330_));
 sky130_fd_sc_hd__and3_1 _12642_ (.A(_05295_),
    .B(_05330_),
    .C(_05271_),
    .X(_05331_));
 sky130_fd_sc_hd__a21oi_1 _12643_ (.A1(_05296_),
    .A2(_05271_),
    .B1(_05330_),
    .Y(_05332_));
 sky130_fd_sc_hd__and3_1 _12644_ (.A(_05295_),
    .B(_05265_),
    .C(_05270_),
    .X(_05333_));
 sky130_fd_sc_hd__a21oi_1 _12645_ (.A1(_05296_),
    .A2(_05265_),
    .B1(_05270_),
    .Y(_05334_));
 sky130_fd_sc_hd__or4_2 _12646_ (.A(_05331_),
    .B(_05332_),
    .C(_05333_),
    .D(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__or2_2 _12647_ (.A(_05233_),
    .B(_05263_),
    .X(_05336_));
 sky130_fd_sc_hd__and2_2 _12648_ (.A(_05227_),
    .B(_05229_),
    .X(_05337_));
 sky130_fd_sc_hd__nor2_1 _12649_ (.A(_05336_),
    .B(_05337_),
    .Y(_05338_));
 sky130_fd_sc_hd__o21ai_4 _12650_ (.A1(_05220_),
    .A2(_05221_),
    .B1(_05223_),
    .Y(_05339_));
 sky130_fd_sc_hd__nand2_2 _12651_ (.A(_05211_),
    .B(_05213_),
    .Y(_05340_));
 sky130_fd_sc_hd__a21oi_2 _12652_ (.A1(_05220_),
    .A2(_05294_),
    .B1(_05280_),
    .Y(_05341_));
 sky130_fd_sc_hd__a31o_1 _12653_ (.A1(_05338_),
    .A2(_05339_),
    .A3(_05340_),
    .B1(_05341_),
    .X(_05342_));
 sky130_fd_sc_hd__xnor2_2 _12654_ (.A(_05218_),
    .B(_05342_),
    .Y(_05343_));
 sky130_fd_sc_hd__inv_2 _12655_ (.A(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__a21o_1 _12656_ (.A1(_05338_),
    .A2(_05339_),
    .B1(_05341_),
    .X(_05345_));
 sky130_fd_sc_hd__xor2_4 _12657_ (.A(_05340_),
    .B(_05345_),
    .X(_05346_));
 sky130_fd_sc_hd__and3b_1 _12658_ (.A_N(_05335_),
    .B(_05344_),
    .C(_05346_),
    .X(_05347_));
 sky130_fd_sc_hd__and4_1 _12659_ (.A(_05310_),
    .B(_05322_),
    .C(_05329_),
    .D(_05347_),
    .X(_05348_));
 sky130_fd_sc_hd__nand2_1 _12660_ (.A(_05305_),
    .B(_05336_),
    .Y(_05349_));
 sky130_fd_sc_hd__xnor2_4 _12661_ (.A(_05337_),
    .B(_05349_),
    .Y(_05350_));
 sky130_fd_sc_hd__or3_1 _12662_ (.A(_05323_),
    .B(_05325_),
    .C(_05327_),
    .X(_05351_));
 sky130_fd_sc_hd__nor2_2 _12663_ (.A(_05341_),
    .B(_05338_),
    .Y(_05352_));
 sky130_fd_sc_hd__xnor2_4 _12664_ (.A(_05339_),
    .B(_05352_),
    .Y(_05353_));
 sky130_fd_sc_hd__or4_1 _12665_ (.A(_05353_),
    .B(_05335_),
    .C(_05343_),
    .D(_05346_),
    .X(_05354_));
 sky130_fd_sc_hd__nor2_1 _12666_ (.A(_05351_),
    .B(_05354_),
    .Y(_05355_));
 sky130_fd_sc_hd__and4_1 _12667_ (.A(_05310_),
    .B(_05322_),
    .C(_05350_),
    .D(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__inv_2 _12668_ (.A(_05346_),
    .Y(_05357_));
 sky130_fd_sc_hd__and4bb_1 _12669_ (.A_N(_05351_),
    .B_N(_05335_),
    .C(_05344_),
    .D(_05357_),
    .X(_05358_));
 sky130_fd_sc_hd__and4_1 _12670_ (.A(_05310_),
    .B(_05322_),
    .C(_05353_),
    .D(_05358_),
    .X(_05359_));
 sky130_fd_sc_hd__nor3_2 _12671_ (.A(_05348_),
    .B(_05356_),
    .C(_05359_),
    .Y(_05360_));
 sky130_fd_sc_hd__nand2_2 _12672_ (.A(_05310_),
    .B(_05322_),
    .Y(_05361_));
 sky130_fd_sc_hd__inv_2 _12673_ (.A(_05350_),
    .Y(_05362_));
 sky130_fd_sc_hd__nand2_2 _12674_ (.A(_05362_),
    .B(_05355_),
    .Y(_05363_));
 sky130_fd_sc_hd__and2_1 _12675_ (.A(_05237_),
    .B(_05239_),
    .X(_05364_));
 sky130_fd_sc_hd__and3_1 _12676_ (.A(_05295_),
    .B(_05364_),
    .C(_05262_),
    .X(_05365_));
 sky130_fd_sc_hd__a21oi_2 _12677_ (.A1(_05296_),
    .A2(_05262_),
    .B1(_05364_),
    .Y(_05366_));
 sky130_fd_sc_hd__and3_1 _12678_ (.A(_05296_),
    .B(_05233_),
    .C(_05263_),
    .X(_05367_));
 sky130_fd_sc_hd__a21oi_1 _12679_ (.A1(_05296_),
    .A2(_05263_),
    .B1(_05233_),
    .Y(_05368_));
 sky130_fd_sc_hd__o22ai_1 _12680_ (.A1(_05365_),
    .A2(_05366_),
    .B1(_05367_),
    .B2(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__a21o_2 _12681_ (.A1(_03790_),
    .A2(_05242_),
    .B1(_05244_),
    .X(_05370_));
 sky130_fd_sc_hd__o21a_1 _12682_ (.A1(_05261_),
    .A2(_05249_),
    .B1(_05295_),
    .X(_05371_));
 sky130_fd_sc_hd__xor2_4 _12683_ (.A(_05370_),
    .B(_05371_),
    .X(_05372_));
 sky130_fd_sc_hd__or2_1 _12684_ (.A(_05369_),
    .B(_05372_),
    .X(_05373_));
 sky130_fd_sc_hd__nand2_1 _12685_ (.A(_05305_),
    .B(_05261_),
    .Y(_05374_));
 sky130_fd_sc_hd__xnor2_4 _12686_ (.A(_05249_),
    .B(_05374_),
    .Y(_05375_));
 sky130_fd_sc_hd__or2_1 _12687_ (.A(_05373_),
    .B(_05375_),
    .X(_05376_));
 sky130_fd_sc_hd__o21ai_2 _12688_ (.A1(_05253_),
    .A2(_05255_),
    .B1(_05305_),
    .Y(_05377_));
 sky130_fd_sc_hd__xnor2_4 _12689_ (.A(_05251_),
    .B(_05377_),
    .Y(_05378_));
 sky130_fd_sc_hd__inv_2 _12690_ (.A(_05378_),
    .Y(_05379_));
 sky130_fd_sc_hd__nand2_1 _12691_ (.A(_05305_),
    .B(_05256_),
    .Y(_05380_));
 sky130_fd_sc_hd__xnor2_4 _12692_ (.A(_05260_),
    .B(_05380_),
    .Y(_05381_));
 sky130_fd_sc_hd__or3_1 _12693_ (.A(_05376_),
    .B(_05379_),
    .C(_05381_),
    .X(_05382_));
 sky130_fd_sc_hd__xnor2_2 _12694_ (.A(_05284_),
    .B(_05316_),
    .Y(_05383_));
 sky130_fd_sc_hd__nand2_1 _12695_ (.A(_05305_),
    .B(_05253_),
    .Y(_05384_));
 sky130_fd_sc_hd__xor2_1 _12696_ (.A(_05255_),
    .B(_05384_),
    .X(_05385_));
 sky130_fd_sc_hd__or3_1 _12697_ (.A(_05378_),
    .B(_05381_),
    .C(_05385_),
    .X(_05386_));
 sky130_fd_sc_hd__or4_1 _12698_ (.A(_05369_),
    .B(_05372_),
    .C(_05350_),
    .D(_05375_),
    .X(_05387_));
 sky130_fd_sc_hd__or4_1 _12699_ (.A(_05351_),
    .B(_05354_),
    .C(_05386_),
    .D(_05387_),
    .X(_05388_));
 sky130_fd_sc_hd__inv_2 _12700_ (.A(_05381_),
    .Y(_05389_));
 sky130_fd_sc_hd__or4_1 _12701_ (.A(_05351_),
    .B(_05354_),
    .C(_05389_),
    .D(_05387_),
    .X(_05390_));
 sky130_fd_sc_hd__nand4_1 _12702_ (.A(_05298_),
    .B(_05300_),
    .C(_05307_),
    .D(_05309_),
    .Y(_05391_));
 sky130_fd_sc_hd__a41o_1 _12703_ (.A1(_05322_),
    .A2(_05383_),
    .A3(_05388_),
    .A4(_05390_),
    .B1(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__o31a_1 _12704_ (.A1(_05361_),
    .A2(_05363_),
    .A3(_05382_),
    .B1(_05392_),
    .X(_05393_));
 sky130_fd_sc_hd__inv_2 _12705_ (.A(_05253_),
    .Y(_05394_));
 sky130_fd_sc_hd__xnor2_1 _12706_ (.A(_05255_),
    .B(_05384_),
    .Y(_05395_));
 sky130_fd_sc_hd__or4_1 _12707_ (.A(_05394_),
    .B(_05378_),
    .C(_05381_),
    .D(_05395_),
    .X(_05396_));
 sky130_fd_sc_hd__or4_2 _12708_ (.A(_05361_),
    .B(_05363_),
    .C(_05376_),
    .D(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__or4_1 _12709_ (.A(_05361_),
    .B(_05351_),
    .C(_05335_),
    .D(_05344_),
    .X(_05398_));
 sky130_fd_sc_hd__and4_1 _12710_ (.A(_05360_),
    .B(_05393_),
    .C(_05397_),
    .D(_05398_),
    .X(_05399_));
 sky130_fd_sc_hd__or3_1 _12711_ (.A(_05336_),
    .B(_05361_),
    .C(_05363_),
    .X(_05400_));
 sky130_fd_sc_hd__buf_4 _12712_ (.A(_05400_),
    .X(_05401_));
 sky130_fd_sc_hd__and2_1 _12713_ (.A(_05310_),
    .B(_05322_),
    .X(_05402_));
 sky130_fd_sc_hd__o211ai_1 _12714_ (.A1(_05328_),
    .A2(_05335_),
    .B1(_05402_),
    .C1(_05383_),
    .Y(_05403_));
 sky130_fd_sc_hd__and4_2 _12715_ (.A(_05360_),
    .B(_05398_),
    .C(_05401_),
    .D(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__nor2_2 _12716_ (.A(_05399_),
    .B(_05404_),
    .Y(_05405_));
 sky130_fd_sc_hd__nand2_2 _12717_ (.A(_05399_),
    .B(_05404_),
    .Y(_05406_));
 sky130_fd_sc_hd__or2b_1 _12718_ (.A(_05405_),
    .B_N(_05406_),
    .X(_05407_));
 sky130_fd_sc_hd__buf_2 _12719_ (.A(_05407_),
    .X(_05408_));
 sky130_fd_sc_hd__or4b_1 _12720_ (.A(_05373_),
    .B(_05361_),
    .C(_05363_),
    .D_N(_05375_),
    .X(_05409_));
 sky130_fd_sc_hd__nand3b_2 _12721_ (.A_N(_05356_),
    .B(_05397_),
    .C(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__nand2_1 _12722_ (.A(_05402_),
    .B(_05323_),
    .Y(_05411_));
 sky130_fd_sc_hd__xor2_1 _12723_ (.A(_05292_),
    .B(_05299_),
    .X(_05412_));
 sky130_fd_sc_hd__nand2_1 _12724_ (.A(_05298_),
    .B(_05412_),
    .Y(_05413_));
 sky130_fd_sc_hd__o311a_1 _12725_ (.A1(_05391_),
    .A2(_05314_),
    .A3(_05318_),
    .B1(_05413_),
    .C1(_05307_),
    .X(_05414_));
 sky130_fd_sc_hd__and3b_1 _12726_ (.A_N(_05348_),
    .B(_05411_),
    .C(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__or2_2 _12727_ (.A(_05361_),
    .B(_05363_),
    .X(_05416_));
 sky130_fd_sc_hd__nor2_4 _12728_ (.A(_05365_),
    .B(_05366_),
    .Y(_05417_));
 sky130_fd_sc_hd__or2_1 _12729_ (.A(_05367_),
    .B(_05368_),
    .X(_05418_));
 sky130_fd_sc_hd__nand2_1 _12730_ (.A(_05417_),
    .B(_05418_),
    .Y(_05419_));
 sky130_fd_sc_hd__inv_2 _12731_ (.A(_05327_),
    .Y(_05420_));
 sky130_fd_sc_hd__or4_1 _12732_ (.A(_05361_),
    .B(_05323_),
    .C(_05325_),
    .D(_05420_),
    .X(_05421_));
 sky130_fd_sc_hd__or2_2 _12733_ (.A(_05331_),
    .B(_05332_),
    .X(_05422_));
 sky130_fd_sc_hd__nor2_1 _12734_ (.A(_05333_),
    .B(_05334_),
    .Y(_05423_));
 sky130_fd_sc_hd__or4_1 _12735_ (.A(_05361_),
    .B(_05351_),
    .C(_05422_),
    .D(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__or3_1 _12736_ (.A(_05361_),
    .B(_05363_),
    .C(_05382_),
    .X(_05425_));
 sky130_fd_sc_hd__o2111a_1 _12737_ (.A1(_05416_),
    .A2(_05419_),
    .B1(_05421_),
    .C1(_05424_),
    .D1(_05425_),
    .X(_05426_));
 sky130_fd_sc_hd__and3b_1 _12738_ (.A_N(_05410_),
    .B(_05415_),
    .C(_05426_),
    .X(_05427_));
 sky130_fd_sc_hd__clkbuf_2 _12739_ (.A(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__clkbuf_4 _12740_ (.A(_05428_),
    .X(_05429_));
 sky130_fd_sc_hd__clkbuf_4 _12741_ (.A(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__buf_2 _12742_ (.A(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__buf_2 _12743_ (.A(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__nor2_2 _12744_ (.A(_05336_),
    .B(_05416_),
    .Y(_05433_));
 sky130_fd_sc_hd__buf_4 _12745_ (.A(_05433_),
    .X(_05434_));
 sky130_fd_sc_hd__xnor2_1 _12746_ (.A(_05315_),
    .B(_05317_),
    .Y(_05435_));
 sky130_fd_sc_hd__or3_1 _12747_ (.A(_05391_),
    .B(_05314_),
    .C(_05435_),
    .X(_05436_));
 sky130_fd_sc_hd__a31oi_2 _12748_ (.A1(_05321_),
    .A2(_05383_),
    .A3(_05388_),
    .B1(_05436_),
    .Y(_05437_));
 sky130_fd_sc_hd__nor2_1 _12749_ (.A(_05367_),
    .B(_05368_),
    .Y(_05438_));
 sky130_fd_sc_hd__nor2_1 _12750_ (.A(_05417_),
    .B(_05438_),
    .Y(_05439_));
 sky130_fd_sc_hd__nor2_2 _12751_ (.A(_05361_),
    .B(_05363_),
    .Y(_05440_));
 sky130_fd_sc_hd__and3_1 _12752_ (.A(_05402_),
    .B(_05329_),
    .C(_05335_),
    .X(_05441_));
 sky130_fd_sc_hd__a21boi_1 _12753_ (.A1(_05298_),
    .A2(_05300_),
    .B1_N(_05307_),
    .Y(_05442_));
 sky130_fd_sc_hd__a311o_1 _12754_ (.A1(_05439_),
    .A2(_05372_),
    .A3(_05440_),
    .B1(_05441_),
    .C1(_05442_),
    .X(_05443_));
 sky130_fd_sc_hd__nor4_4 _12755_ (.A(_05359_),
    .B(_05410_),
    .C(_05437_),
    .D(_05443_),
    .Y(_05444_));
 sky130_fd_sc_hd__a21o_1 _12756_ (.A1(_05444_),
    .A2(_05428_),
    .B1(_05399_),
    .X(_05445_));
 sky130_fd_sc_hd__and2_1 _12757_ (.A(_05404_),
    .B(_05445_),
    .X(_05446_));
 sky130_fd_sc_hd__buf_4 _12758_ (.A(_05446_),
    .X(_05447_));
 sky130_fd_sc_hd__clkbuf_4 _12759_ (.A(_05428_),
    .X(_05448_));
 sky130_fd_sc_hd__mux2_1 _12760_ (.A0(_05346_),
    .A1(_05353_),
    .S(_05448_),
    .X(_05449_));
 sky130_fd_sc_hd__or2_1 _12761_ (.A(_05333_),
    .B(_05334_),
    .X(_05450_));
 sky130_fd_sc_hd__mux2_1 _12762_ (.A0(_05450_),
    .A1(_05343_),
    .S(_05448_),
    .X(_05451_));
 sky130_fd_sc_hd__or4_2 _12763_ (.A(_05359_),
    .B(_05410_),
    .C(_05437_),
    .D(_05443_),
    .X(_05452_));
 sky130_fd_sc_hd__xnor2_2 _12764_ (.A(_05452_),
    .B(_05428_),
    .Y(_05453_));
 sky130_fd_sc_hd__mux2_1 _12765_ (.A0(_05449_),
    .A1(_05451_),
    .S(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__mux2_1 _12766_ (.A0(_05327_),
    .A1(_05422_),
    .S(_05448_),
    .X(_05455_));
 sky130_fd_sc_hd__mux2_1 _12767_ (.A0(_05323_),
    .A1(_05325_),
    .S(_05448_),
    .X(_05456_));
 sky130_fd_sc_hd__mux2_1 _12768_ (.A0(_05455_),
    .A1(_05456_),
    .S(_05453_),
    .X(_05457_));
 sky130_fd_sc_hd__nand4_2 _12769_ (.A(_05360_),
    .B(_05393_),
    .C(_05397_),
    .D(_05398_),
    .Y(_05458_));
 sky130_fd_sc_hd__or3b_2 _12770_ (.A(_05458_),
    .B(_05452_),
    .C_N(_05428_),
    .X(_05459_));
 sky130_fd_sc_hd__nand2_1 _12771_ (.A(_05459_),
    .B(_05445_),
    .Y(_05460_));
 sky130_fd_sc_hd__mux2_1 _12772_ (.A0(_05454_),
    .A1(_05457_),
    .S(_05460_),
    .X(_05461_));
 sky130_fd_sc_hd__clkbuf_4 _12773_ (.A(_05452_),
    .X(_05462_));
 sky130_fd_sc_hd__clkbuf_4 _12774_ (.A(_05448_),
    .X(_05463_));
 sky130_fd_sc_hd__mux4_1 _12775_ (.A0(_05375_),
    .A1(_05378_),
    .A2(_05395_),
    .A3(_05381_),
    .S0(_05462_),
    .S1(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__mux4_1 _12776_ (.A0(_05417_),
    .A1(_05438_),
    .A2(_05350_),
    .A3(_05372_),
    .S0(_05448_),
    .S1(_05444_),
    .X(_05465_));
 sky130_fd_sc_hd__a21o_1 _12777_ (.A1(_05459_),
    .A2(_05445_),
    .B1(_05465_),
    .X(_05466_));
 sky130_fd_sc_hd__nand2_1 _12778_ (.A(_05404_),
    .B(_05445_),
    .Y(_05467_));
 sky130_fd_sc_hd__o211a_1 _12779_ (.A1(_05460_),
    .A2(_05464_),
    .B1(_05466_),
    .C1(_05467_),
    .X(_05468_));
 sky130_fd_sc_hd__or3_1 _12780_ (.A(_05348_),
    .B(_05356_),
    .C(_05359_),
    .X(_05469_));
 sky130_fd_sc_hd__clkbuf_4 _12781_ (.A(_05469_),
    .X(_05470_));
 sky130_fd_sc_hd__a211o_2 _12782_ (.A1(_05447_),
    .A2(_05461_),
    .B1(_05468_),
    .C1(_05470_),
    .X(_05471_));
 sky130_fd_sc_hd__mux2_1 _12783_ (.A0(_05394_),
    .A1(_05385_),
    .S(_05429_),
    .X(_05472_));
 sky130_fd_sc_hd__nor2_1 _12784_ (.A(_05462_),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__or2_2 _12785_ (.A(_05360_),
    .B(_05473_),
    .X(_05474_));
 sky130_fd_sc_hd__mux4_1 _12786_ (.A0(_05438_),
    .A1(_05372_),
    .A2(_05375_),
    .A3(_05417_),
    .S0(_05462_),
    .S1(_05463_),
    .X(_05475_));
 sky130_fd_sc_hd__mux4_1 _12787_ (.A0(_05381_),
    .A1(_05395_),
    .A2(_05253_),
    .A3(_05378_),
    .S0(_05462_),
    .S1(_05463_),
    .X(_05476_));
 sky130_fd_sc_hd__and2_1 _12788_ (.A(_05459_),
    .B(_05445_),
    .X(_05477_));
 sky130_fd_sc_hd__buf_2 _12789_ (.A(_05477_),
    .X(_05478_));
 sky130_fd_sc_hd__mux2_1 _12790_ (.A0(_05475_),
    .A1(_05476_),
    .S(_05478_),
    .X(_05479_));
 sky130_fd_sc_hd__nand2_2 _12791_ (.A(_05416_),
    .B(_05360_),
    .Y(_05480_));
 sky130_fd_sc_hd__a21o_1 _12792_ (.A1(_05404_),
    .A2(_05445_),
    .B1(_05470_),
    .X(_05481_));
 sky130_fd_sc_hd__nor2_1 _12793_ (.A(_05480_),
    .B(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__mux4_1 _12794_ (.A0(_05353_),
    .A1(_05343_),
    .A2(_05346_),
    .A3(_05350_),
    .S0(_05444_),
    .S1(_05463_),
    .X(_05483_));
 sky130_fd_sc_hd__mux2_1 _12795_ (.A0(_05422_),
    .A1(_05450_),
    .S(_05448_),
    .X(_05484_));
 sky130_fd_sc_hd__mux2_1 _12796_ (.A0(_05325_),
    .A1(_05327_),
    .S(_05448_),
    .X(_05485_));
 sky130_fd_sc_hd__mux2_1 _12797_ (.A0(_05484_),
    .A1(_05485_),
    .S(_05453_),
    .X(_05486_));
 sky130_fd_sc_hd__mux2_2 _12798_ (.A0(_05483_),
    .A1(_05486_),
    .S(_05460_),
    .X(_05487_));
 sky130_fd_sc_hd__o22a_2 _12799_ (.A1(_05447_),
    .A2(_05479_),
    .B1(_05482_),
    .B2(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__a21o_2 _12800_ (.A1(_05471_),
    .A2(_05474_),
    .B1(_05488_),
    .X(_05489_));
 sky130_fd_sc_hd__mux2_1 _12801_ (.A0(_05344_),
    .A1(_05357_),
    .S(_05429_),
    .X(_05490_));
 sky130_fd_sc_hd__clkinv_2 _12802_ (.A(_05422_),
    .Y(_05491_));
 sky130_fd_sc_hd__mux2_1 _12803_ (.A0(_05491_),
    .A1(_05423_),
    .S(_05429_),
    .X(_05492_));
 sky130_fd_sc_hd__mux2_1 _12804_ (.A0(_05490_),
    .A1(_05492_),
    .S(_05453_),
    .X(_05493_));
 sky130_fd_sc_hd__clkinv_2 _12805_ (.A(_05325_),
    .Y(_05494_));
 sky130_fd_sc_hd__mux2_1 _12806_ (.A0(_05494_),
    .A1(_05420_),
    .S(_05429_),
    .X(_05495_));
 sky130_fd_sc_hd__mux2_1 _12807_ (.A0(_05321_),
    .A1(_05383_),
    .S(_05429_),
    .X(_05496_));
 sky130_fd_sc_hd__buf_2 _12808_ (.A(_05453_),
    .X(_05497_));
 sky130_fd_sc_hd__mux2_1 _12809_ (.A0(_05495_),
    .A1(_05496_),
    .S(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__buf_2 _12810_ (.A(_05460_),
    .X(_05499_));
 sky130_fd_sc_hd__mux2_1 _12811_ (.A0(_05493_),
    .A1(_05498_),
    .S(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__buf_2 _12812_ (.A(_05444_),
    .X(_05501_));
 sky130_fd_sc_hd__mux2_1 _12813_ (.A0(_05395_),
    .A1(_05378_),
    .S(_05429_),
    .X(_05502_));
 sky130_fd_sc_hd__and3_1 _12814_ (.A(_05253_),
    .B(_05462_),
    .C(_05463_),
    .X(_05503_));
 sky130_fd_sc_hd__a21oi_1 _12815_ (.A1(_05501_),
    .A2(_05502_),
    .B1(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__inv_2 _12816_ (.A(_05353_),
    .Y(_05505_));
 sky130_fd_sc_hd__inv_2 _12817_ (.A(_05417_),
    .Y(_05506_));
 sky130_fd_sc_hd__mux4_1 _12818_ (.A0(_05418_),
    .A1(_05362_),
    .A2(_05505_),
    .A3(_05506_),
    .S0(_05429_),
    .S1(_05444_),
    .X(_05507_));
 sky130_fd_sc_hd__mux4_1 _12819_ (.A0(_05372_),
    .A1(_05378_),
    .A2(_05381_),
    .A3(_05375_),
    .S0(_05428_),
    .S1(_05452_),
    .X(_05508_));
 sky130_fd_sc_hd__inv_2 _12820_ (.A(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hd__mux2_1 _12821_ (.A0(_05507_),
    .A1(_05509_),
    .S(_05478_),
    .X(_05510_));
 sky130_fd_sc_hd__o22a_1 _12822_ (.A1(_05360_),
    .A2(_05504_),
    .B1(_05510_),
    .B2(_05481_),
    .X(_05511_));
 sky130_fd_sc_hd__o21ai_1 _12823_ (.A1(_05467_),
    .A2(_05500_),
    .B1(_05511_),
    .Y(_05512_));
 sky130_fd_sc_hd__mux2_1 _12824_ (.A0(_05379_),
    .A1(_05389_),
    .S(_05463_),
    .X(_05513_));
 sky130_fd_sc_hd__mux2_2 _12825_ (.A0(_05513_),
    .A1(_05472_),
    .S(_05462_),
    .X(_05514_));
 sky130_fd_sc_hd__nand2_1 _12826_ (.A(_05444_),
    .B(_05463_),
    .Y(_05515_));
 sky130_fd_sc_hd__or2_1 _12827_ (.A(_05444_),
    .B(_05429_),
    .X(_05516_));
 sky130_fd_sc_hd__nand2_2 _12828_ (.A(_05515_),
    .B(_05516_),
    .Y(_05517_));
 sky130_fd_sc_hd__nand2_1 _12829_ (.A(_05497_),
    .B(_05455_),
    .Y(_05518_));
 sky130_fd_sc_hd__a21boi_1 _12830_ (.A1(_05517_),
    .A2(_05451_),
    .B1_N(_05518_),
    .Y(_05519_));
 sky130_fd_sc_hd__or2_1 _12831_ (.A(_05499_),
    .B(_05519_),
    .X(_05520_));
 sky130_fd_sc_hd__mux4_1 _12832_ (.A0(_05350_),
    .A1(_05353_),
    .A2(_05346_),
    .A3(_05438_),
    .S0(_05429_),
    .S1(_05501_),
    .X(_05521_));
 sky130_fd_sc_hd__mux4_1 _12833_ (.A0(_05417_),
    .A1(_05375_),
    .A2(_05381_),
    .A3(_05372_),
    .S0(_05462_),
    .S1(_05430_),
    .X(_05522_));
 sky130_fd_sc_hd__mux2_1 _12834_ (.A0(_05521_),
    .A1(_05522_),
    .S(_05478_),
    .X(_05523_));
 sky130_fd_sc_hd__nor2_1 _12835_ (.A(_05447_),
    .B(_05523_),
    .Y(_05524_));
 sky130_fd_sc_hd__a221oi_4 _12836_ (.A1(_05470_),
    .A2(_05514_),
    .B1(_05520_),
    .B2(_05447_),
    .C1(_05524_),
    .Y(_05525_));
 sky130_fd_sc_hd__a21o_2 _12837_ (.A1(_05489_),
    .A2(_05512_),
    .B1(_05525_),
    .X(_05526_));
 sky130_fd_sc_hd__clkbuf_4 _12838_ (.A(_05478_),
    .X(_05527_));
 sky130_fd_sc_hd__mux2_1 _12839_ (.A0(_05378_),
    .A1(_05381_),
    .S(_05448_),
    .X(_05528_));
 sky130_fd_sc_hd__mux2_1 _12840_ (.A0(_05375_),
    .A1(_05372_),
    .S(_05448_),
    .X(_05529_));
 sky130_fd_sc_hd__mux2_1 _12841_ (.A0(_05528_),
    .A1(_05529_),
    .S(_05444_),
    .X(_05530_));
 sky130_fd_sc_hd__buf_2 _12842_ (.A(_05399_),
    .X(_05531_));
 sky130_fd_sc_hd__mux2_1 _12843_ (.A0(_05530_),
    .A1(_05473_),
    .S(_05531_),
    .X(_05532_));
 sky130_fd_sc_hd__and2_1 _12844_ (.A(_05480_),
    .B(_05532_),
    .X(_05533_));
 sky130_fd_sc_hd__or2_1 _12845_ (.A(_05478_),
    .B(_05454_),
    .X(_05534_));
 sky130_fd_sc_hd__nor2_2 _12846_ (.A(_05470_),
    .B(_05447_),
    .Y(_05535_));
 sky130_fd_sc_hd__o211a_1 _12847_ (.A1(_05499_),
    .A2(_05465_),
    .B1(_05534_),
    .C1(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__a211oi_4 _12848_ (.A1(_05527_),
    .A2(_05457_),
    .B1(_05533_),
    .C1(_05536_),
    .Y(_05537_));
 sky130_fd_sc_hd__nor2_2 _12849_ (.A(_05440_),
    .B(_05470_),
    .Y(_05538_));
 sky130_fd_sc_hd__mux2_1 _12850_ (.A0(_05381_),
    .A1(_05375_),
    .S(_05463_),
    .X(_05539_));
 sky130_fd_sc_hd__mux2_1 _12851_ (.A0(_05539_),
    .A1(_05502_),
    .S(_05462_),
    .X(_05540_));
 sky130_fd_sc_hd__o2bb2a_1 _12852_ (.A1_N(_05458_),
    .A2_N(_05540_),
    .B1(_05459_),
    .B2(_05394_),
    .X(_05541_));
 sky130_fd_sc_hd__mux2_1 _12853_ (.A0(_05483_),
    .A1(_05475_),
    .S(_05478_),
    .X(_05542_));
 sky130_fd_sc_hd__a22o_1 _12854_ (.A1(_05527_),
    .A2(_05486_),
    .B1(_05467_),
    .B2(_05538_),
    .X(_05543_));
 sky130_fd_sc_hd__o21ai_1 _12855_ (.A1(_05481_),
    .A2(_05542_),
    .B1(_05543_),
    .Y(_05544_));
 sky130_fd_sc_hd__o21a_2 _12856_ (.A1(_05538_),
    .A2(_05541_),
    .B1(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__nor2_1 _12857_ (.A(_05537_),
    .B(_05545_),
    .Y(_05546_));
 sky130_fd_sc_hd__mux2_1 _12858_ (.A0(_05372_),
    .A1(_05417_),
    .S(_05463_),
    .X(_05547_));
 sky130_fd_sc_hd__mux2_1 _12859_ (.A0(_05539_),
    .A1(_05547_),
    .S(_05501_),
    .X(_05548_));
 sky130_fd_sc_hd__o2bb2a_1 _12860_ (.A1_N(_05405_),
    .A2_N(_05548_),
    .B1(_05504_),
    .B2(_05406_),
    .X(_05549_));
 sky130_fd_sc_hd__mux2_1 _12861_ (.A0(_05493_),
    .A1(_05507_),
    .S(_05478_),
    .X(_05550_));
 sky130_fd_sc_hd__or2_1 _12862_ (.A(_05481_),
    .B(_05550_),
    .X(_05551_));
 sky130_fd_sc_hd__o221a_1 _12863_ (.A1(_05499_),
    .A2(_05498_),
    .B1(_05549_),
    .B2(_05538_),
    .C1(_05551_),
    .X(_05552_));
 sky130_fd_sc_hd__clkinv_2 _12864_ (.A(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__mux2_1 _12865_ (.A0(_05318_),
    .A1(_05321_),
    .S(_05430_),
    .X(_05554_));
 sky130_fd_sc_hd__nor2_1 _12866_ (.A(_05497_),
    .B(_05456_),
    .Y(_05555_));
 sky130_fd_sc_hd__a21o_1 _12867_ (.A1(_05497_),
    .A2(_05554_),
    .B1(_05555_),
    .X(_05556_));
 sky130_fd_sc_hd__nor2_1 _12868_ (.A(_05499_),
    .B(_05521_),
    .Y(_05557_));
 sky130_fd_sc_hd__a211o_1 _12869_ (.A1(_05499_),
    .A2(_05519_),
    .B1(_05557_),
    .C1(_05481_),
    .X(_05558_));
 sky130_fd_sc_hd__nor2_1 _12870_ (.A(_05406_),
    .B(_05514_),
    .Y(_05559_));
 sky130_fd_sc_hd__mux2_1 _12871_ (.A0(_05506_),
    .A1(_05418_),
    .S(_05430_),
    .X(_05560_));
 sky130_fd_sc_hd__nand2_1 _12872_ (.A(_05501_),
    .B(_05560_),
    .Y(_05561_));
 sky130_fd_sc_hd__o211a_1 _12873_ (.A1(_05501_),
    .A2(_05529_),
    .B1(_05561_),
    .C1(_05405_),
    .X(_05562_));
 sky130_fd_sc_hd__o21ai_1 _12874_ (.A1(_05559_),
    .A2(_05562_),
    .B1(_05480_),
    .Y(_05563_));
 sky130_fd_sc_hd__o211a_2 _12875_ (.A1(_05556_),
    .A2(_05499_),
    .B1(_05558_),
    .C1(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__inv_2 _12876_ (.A(_05564_),
    .Y(_05565_));
 sky130_fd_sc_hd__a31o_1 _12877_ (.A1(_05526_),
    .A2(_05546_),
    .A3(_05553_),
    .B1(_05565_),
    .X(_05566_));
 sky130_fd_sc_hd__buf_2 _12878_ (.A(_05566_),
    .X(_05567_));
 sky130_fd_sc_hd__nor2_2 _12879_ (.A(_05440_),
    .B(_05405_),
    .Y(_05568_));
 sky130_fd_sc_hd__nor2b_1 _12880_ (.A(_05405_),
    .B_N(_05406_),
    .Y(_05569_));
 sky130_fd_sc_hd__o21a_1 _12881_ (.A1(_05531_),
    .A2(_05504_),
    .B1(_05569_),
    .X(_05570_));
 sky130_fd_sc_hd__mux2_1 _12882_ (.A0(_05418_),
    .A1(_05362_),
    .S(_05463_),
    .X(_05571_));
 sky130_fd_sc_hd__nor2_1 _12883_ (.A(_05353_),
    .B(_05430_),
    .Y(_05572_));
 sky130_fd_sc_hd__a211o_1 _12884_ (.A1(_05357_),
    .A2(_05430_),
    .B1(_05572_),
    .C1(_05462_),
    .X(_05573_));
 sky130_fd_sc_hd__o211a_1 _12885_ (.A1(_05501_),
    .A2(_05571_),
    .B1(_05573_),
    .C1(_05405_),
    .X(_05574_));
 sky130_fd_sc_hd__nor2_1 _12886_ (.A(_05406_),
    .B(_05548_),
    .Y(_05575_));
 sky130_fd_sc_hd__or4_1 _12887_ (.A(_05568_),
    .B(_05570_),
    .C(_05574_),
    .D(_05575_),
    .X(_05576_));
 sky130_fd_sc_hd__buf_2 _12888_ (.A(_05481_),
    .X(_05577_));
 sky130_fd_sc_hd__mux2_1 _12889_ (.A0(_05314_),
    .A1(_05435_),
    .S(_05430_),
    .X(_05578_));
 sky130_fd_sc_hd__nand2_1 _12890_ (.A(_05517_),
    .B(_05578_),
    .Y(_05579_));
 sky130_fd_sc_hd__mux2_1 _12891_ (.A0(_05298_),
    .A1(_05300_),
    .S(_05430_),
    .X(_05580_));
 sky130_fd_sc_hd__o211a_1 _12892_ (.A1(_05577_),
    .A2(_05500_),
    .B1(_05579_),
    .C1(_05580_),
    .X(_05581_));
 sky130_fd_sc_hd__mux2_1 _12893_ (.A0(_05576_),
    .A1(_05581_),
    .S(_05538_),
    .X(_05582_));
 sky130_fd_sc_hd__inv_2 _12894_ (.A(_05582_),
    .Y(_05583_));
 sky130_fd_sc_hd__nor2_1 _12895_ (.A(_05497_),
    .B(_05496_),
    .Y(_05584_));
 sky130_fd_sc_hd__a221o_1 _12896_ (.A1(_05487_),
    .A2(_05535_),
    .B1(_05578_),
    .B2(_05497_),
    .C1(_05584_),
    .X(_05585_));
 sky130_fd_sc_hd__clkbuf_4 _12897_ (.A(_05462_),
    .X(_05586_));
 sky130_fd_sc_hd__o21ai_1 _12898_ (.A1(_05586_),
    .A2(_05571_),
    .B1(_05405_),
    .Y(_05587_));
 sky130_fd_sc_hd__a21o_1 _12899_ (.A1(_05586_),
    .A2(_05547_),
    .B1(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__a41o_1 _12900_ (.A1(_05253_),
    .A2(_05458_),
    .A3(_05501_),
    .A4(_05431_),
    .B1(_05407_),
    .X(_05589_));
 sky130_fd_sc_hd__o2111a_1 _12901_ (.A1(_05406_),
    .A2(_05540_),
    .B1(_05588_),
    .C1(_05589_),
    .D1(_05480_),
    .X(_05590_));
 sky130_fd_sc_hd__nor2_2 _12902_ (.A(_05585_),
    .B(_05590_),
    .Y(_05591_));
 sky130_fd_sc_hd__nand2_1 _12903_ (.A(_05535_),
    .B(_05461_),
    .Y(_05592_));
 sky130_fd_sc_hd__inv_2 _12904_ (.A(_05431_),
    .Y(_05593_));
 sky130_fd_sc_hd__nor2_1 _12905_ (.A(_05314_),
    .B(_05593_),
    .Y(_05594_));
 sky130_fd_sc_hd__o21ai_1 _12906_ (.A1(_05412_),
    .A2(_05431_),
    .B1(_05497_),
    .Y(_05595_));
 sky130_fd_sc_hd__o22a_1 _12907_ (.A1(_05497_),
    .A2(_05554_),
    .B1(_05594_),
    .B2(_05595_),
    .X(_05596_));
 sky130_fd_sc_hd__o31ai_1 _12908_ (.A1(_05531_),
    .A2(_05586_),
    .A3(_05472_),
    .B1(_05569_),
    .Y(_05597_));
 sky130_fd_sc_hd__o21ai_1 _12909_ (.A1(_05406_),
    .A2(_05530_),
    .B1(_05597_),
    .Y(_05598_));
 sky130_fd_sc_hd__nor2_1 _12910_ (.A(_05350_),
    .B(_05430_),
    .Y(_05599_));
 sky130_fd_sc_hd__a211o_1 _12911_ (.A1(_05505_),
    .A2(_05430_),
    .B1(_05599_),
    .C1(_05586_),
    .X(_05600_));
 sky130_fd_sc_hd__o211a_1 _12912_ (.A1(_05501_),
    .A2(_05560_),
    .B1(_05600_),
    .C1(_05405_),
    .X(_05601_));
 sky130_fd_sc_hd__clkbuf_2 _12913_ (.A(_05480_),
    .X(_05602_));
 sky130_fd_sc_hd__o31a_1 _12914_ (.A1(_05568_),
    .A2(_05598_),
    .A3(_05601_),
    .B1(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__a31o_2 _12915_ (.A1(_05538_),
    .A2(_05592_),
    .A3(_05596_),
    .B1(_05603_),
    .X(_05604_));
 sky130_fd_sc_hd__nor2_1 _12916_ (.A(_05591_),
    .B(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hd__and3_1 _12917_ (.A(_05567_),
    .B(_05583_),
    .C(_05605_),
    .X(_05606_));
 sky130_fd_sc_hd__buf_2 _12918_ (.A(_05537_),
    .X(_05607_));
 sky130_fd_sc_hd__clkbuf_4 _12919_ (.A(_05591_),
    .X(_05608_));
 sky130_fd_sc_hd__xnor2_1 _12920_ (.A(_05608_),
    .B(_05566_),
    .Y(_05609_));
 sky130_fd_sc_hd__clkbuf_4 _12921_ (.A(_05609_),
    .X(_05610_));
 sky130_fd_sc_hd__buf_2 _12922_ (.A(_05564_),
    .X(_05611_));
 sky130_fd_sc_hd__clkbuf_4 _12923_ (.A(_05512_),
    .X(_05612_));
 sky130_fd_sc_hd__a21oi_4 _12924_ (.A1(_05489_),
    .A2(_05612_),
    .B1(_05525_),
    .Y(_05613_));
 sky130_fd_sc_hd__or2_1 _12925_ (.A(_05537_),
    .B(_05545_),
    .X(_05614_));
 sky130_fd_sc_hd__nor2_2 _12926_ (.A(_05613_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__clkbuf_4 _12927_ (.A(_05552_),
    .X(_05616_));
 sky130_fd_sc_hd__or3_1 _12928_ (.A(_05613_),
    .B(_05614_),
    .C(_05616_),
    .X(_05617_));
 sky130_fd_sc_hd__buf_2 _12929_ (.A(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__o21a_1 _12930_ (.A1(_05611_),
    .A2(_05615_),
    .B1(_05618_),
    .X(_05619_));
 sky130_fd_sc_hd__or3_1 _12931_ (.A(_05607_),
    .B(_05610_),
    .C(_05619_),
    .X(_05620_));
 sky130_fd_sc_hd__clkbuf_4 _12932_ (.A(_05604_),
    .X(_05621_));
 sky130_fd_sc_hd__xnor2_4 _12933_ (.A(_05526_),
    .B(_05545_),
    .Y(_05622_));
 sky130_fd_sc_hd__or2_1 _12934_ (.A(_05621_),
    .B(_05622_),
    .X(_05623_));
 sky130_fd_sc_hd__clkbuf_4 _12935_ (.A(_05582_),
    .X(_05624_));
 sky130_fd_sc_hd__a221o_4 _12936_ (.A1(_05470_),
    .A2(_05514_),
    .B1(_05520_),
    .B2(_05447_),
    .C1(_05524_),
    .X(_05625_));
 sky130_fd_sc_hd__a21o_1 _12937_ (.A1(_05489_),
    .A2(_05612_),
    .B1(_05625_),
    .X(_05626_));
 sky130_fd_sc_hd__a21oi_4 _12938_ (.A1(_05471_),
    .A2(_05474_),
    .B1(_05488_),
    .Y(_05627_));
 sky130_fd_sc_hd__o21a_1 _12939_ (.A1(_05467_),
    .A2(_05500_),
    .B1(_05511_),
    .X(_05628_));
 sky130_fd_sc_hd__buf_2 _12940_ (.A(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__or3_2 _12941_ (.A(_05627_),
    .B(_05629_),
    .C(_05525_),
    .X(_05630_));
 sky130_fd_sc_hd__and2_1 _12942_ (.A(_05626_),
    .B(_05630_),
    .X(_05631_));
 sky130_fd_sc_hd__nor2_1 _12943_ (.A(_05624_),
    .B(_05631_),
    .Y(_05632_));
 sky130_fd_sc_hd__xnor2_1 _12944_ (.A(_05623_),
    .B(_05632_),
    .Y(_05633_));
 sky130_fd_sc_hd__nand2_4 _12945_ (.A(_05526_),
    .B(_05546_),
    .Y(_05634_));
 sky130_fd_sc_hd__clkbuf_4 _12946_ (.A(_05545_),
    .X(_05635_));
 sky130_fd_sc_hd__o21ai_4 _12947_ (.A1(_05613_),
    .A2(_05635_),
    .B1(_05537_),
    .Y(_05636_));
 sky130_fd_sc_hd__and2_1 _12948_ (.A(_05634_),
    .B(_05636_),
    .X(_05637_));
 sky130_fd_sc_hd__buf_2 _12949_ (.A(_05637_),
    .X(_05638_));
 sky130_fd_sc_hd__nor2_1 _12950_ (.A(_05608_),
    .B(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__xnor2_1 _12951_ (.A(_05613_),
    .B(_05545_),
    .Y(_05640_));
 sky130_fd_sc_hd__clkbuf_4 _12952_ (.A(_05640_),
    .X(_05641_));
 sky130_fd_sc_hd__nand2_1 _12953_ (.A(_05641_),
    .B(_05632_),
    .Y(_05642_));
 sky130_fd_sc_hd__nor2_1 _12954_ (.A(_05621_),
    .B(_05642_),
    .Y(_05643_));
 sky130_fd_sc_hd__a21o_1 _12955_ (.A1(_05633_),
    .A2(_05639_),
    .B1(_05643_),
    .X(_05644_));
 sky130_fd_sc_hd__clkinv_2 _12956_ (.A(_05608_),
    .Y(_05645_));
 sky130_fd_sc_hd__nand2_1 _12957_ (.A(_05611_),
    .B(_05616_),
    .Y(_05646_));
 sky130_fd_sc_hd__a22oi_1 _12958_ (.A1(_05645_),
    .A2(_05634_),
    .B1(_05618_),
    .B2(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__a31o_1 _12959_ (.A1(_05645_),
    .A2(_05634_),
    .A3(_05646_),
    .B1(_05647_),
    .X(_05648_));
 sky130_fd_sc_hd__xnor2_1 _12960_ (.A(_05644_),
    .B(_05648_),
    .Y(_05649_));
 sky130_fd_sc_hd__xnor2_1 _12961_ (.A(_05620_),
    .B(_05649_),
    .Y(_05650_));
 sky130_fd_sc_hd__nand2_2 _12962_ (.A(_05626_),
    .B(_05630_),
    .Y(_05651_));
 sky130_fd_sc_hd__nor2_1 _12963_ (.A(_05624_),
    .B(_05622_),
    .Y(_05652_));
 sky130_fd_sc_hd__or2_1 _12964_ (.A(_05651_),
    .B(_05652_),
    .X(_05653_));
 sky130_fd_sc_hd__nand2_1 _12965_ (.A(_05642_),
    .B(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__nor2_1 _12966_ (.A(_05621_),
    .B(_05638_),
    .Y(_05655_));
 sky130_fd_sc_hd__xor2_1 _12967_ (.A(_05654_),
    .B(_05655_),
    .X(_05656_));
 sky130_fd_sc_hd__and3_2 _12968_ (.A(_05488_),
    .B(_05471_),
    .C(_05474_),
    .X(_05657_));
 sky130_fd_sc_hd__or3_2 _12969_ (.A(_05627_),
    .B(_05582_),
    .C(_05657_),
    .X(_05658_));
 sky130_fd_sc_hd__xnor2_1 _12970_ (.A(_05489_),
    .B(_05628_),
    .Y(_05659_));
 sky130_fd_sc_hd__clkbuf_4 _12971_ (.A(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__xnor2_1 _12972_ (.A(_05633_),
    .B(_05639_),
    .Y(_05661_));
 sky130_fd_sc_hd__or2_1 _12973_ (.A(_05433_),
    .B(_05660_),
    .X(_05662_));
 sky130_fd_sc_hd__or2b_1 _12974_ (.A(_05662_),
    .B_N(_05658_),
    .X(_05663_));
 sky130_fd_sc_hd__o22ai_1 _12975_ (.A1(_05658_),
    .A2(_05660_),
    .B1(_05661_),
    .B2(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__xnor2_1 _12976_ (.A(_05656_),
    .B(_05664_),
    .Y(_05665_));
 sky130_fd_sc_hd__xnor2_1 _12977_ (.A(_05650_),
    .B(_05665_),
    .Y(_05666_));
 sky130_fd_sc_hd__xor2_1 _12978_ (.A(_05661_),
    .B(_05663_),
    .X(_05667_));
 sky130_fd_sc_hd__nor2_4 _12979_ (.A(_05627_),
    .B(_05657_),
    .Y(_05668_));
 sky130_fd_sc_hd__nor2_1 _12980_ (.A(_05624_),
    .B(_05660_),
    .Y(_05669_));
 sky130_fd_sc_hd__xnor2_1 _12981_ (.A(_05668_),
    .B(_05669_),
    .Y(_05670_));
 sky130_fd_sc_hd__nand2_4 _12982_ (.A(_05471_),
    .B(_05474_),
    .Y(_05671_));
 sky130_fd_sc_hd__o22ai_4 _12983_ (.A1(_05447_),
    .A2(_05479_),
    .B1(_05482_),
    .B2(_05487_),
    .Y(_05672_));
 sky130_fd_sc_hd__nor2_1 _12984_ (.A(_05672_),
    .B(_05624_),
    .Y(_05673_));
 sky130_fd_sc_hd__nor2_1 _12985_ (.A(_05604_),
    .B(_05659_),
    .Y(_05674_));
 sky130_fd_sc_hd__xnor2_1 _12986_ (.A(_05488_),
    .B(_05658_),
    .Y(_05675_));
 sky130_fd_sc_hd__a22o_1 _12987_ (.A1(_05671_),
    .A2(_05673_),
    .B1(_05674_),
    .B2(_05675_),
    .X(_05676_));
 sky130_fd_sc_hd__and2b_1 _12988_ (.A_N(_05670_),
    .B(_05676_),
    .X(_05677_));
 sky130_fd_sc_hd__a2bb2o_1 _12989_ (.A1_N(_05621_),
    .A2_N(_05631_),
    .B1(_05641_),
    .B2(_05645_),
    .X(_05678_));
 sky130_fd_sc_hd__a21oi_1 _12990_ (.A1(_05626_),
    .A2(_05630_),
    .B1(_05591_),
    .Y(_05679_));
 sky130_fd_sc_hd__or3b_1 _12991_ (.A(_05604_),
    .B(_05622_),
    .C_N(_05679_),
    .X(_05680_));
 sky130_fd_sc_hd__a21oi_1 _12992_ (.A1(_05634_),
    .A2(_05636_),
    .B1(_05611_),
    .Y(_05681_));
 sky130_fd_sc_hd__nand3_1 _12993_ (.A(_05678_),
    .B(_05680_),
    .C(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__a21o_1 _12994_ (.A1(_05678_),
    .A2(_05680_),
    .B1(_05681_),
    .X(_05683_));
 sky130_fd_sc_hd__xnor2_1 _12995_ (.A(_05670_),
    .B(_05676_),
    .Y(_05684_));
 sky130_fd_sc_hd__and3_1 _12996_ (.A(_05682_),
    .B(_05683_),
    .C(_05684_),
    .X(_05685_));
 sky130_fd_sc_hd__or2_1 _12997_ (.A(_05677_),
    .B(_05685_),
    .X(_05686_));
 sky130_fd_sc_hd__xor2_1 _12998_ (.A(_05667_),
    .B(_05686_),
    .X(_05687_));
 sky130_fd_sc_hd__nand2_1 _12999_ (.A(_05680_),
    .B(_05682_),
    .Y(_05688_));
 sky130_fd_sc_hd__o21ai_1 _13000_ (.A1(_05607_),
    .A2(_05610_),
    .B1(_05619_),
    .Y(_05689_));
 sky130_fd_sc_hd__and2_1 _13001_ (.A(_05620_),
    .B(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__xnor2_1 _13002_ (.A(_05688_),
    .B(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hd__buf_2 _13003_ (.A(_05565_),
    .X(_05692_));
 sky130_fd_sc_hd__or4_1 _13004_ (.A(_05608_),
    .B(_05611_),
    .C(_05537_),
    .D(_05635_),
    .X(_05693_));
 sky130_fd_sc_hd__o21ai_1 _13005_ (.A1(_05692_),
    .A2(_05618_),
    .B1(_05693_),
    .Y(_05694_));
 sky130_fd_sc_hd__xnor2_1 _13006_ (.A(_05691_),
    .B(_05694_),
    .Y(_05695_));
 sky130_fd_sc_hd__and2_1 _13007_ (.A(_05667_),
    .B(_05686_),
    .X(_05696_));
 sky130_fd_sc_hd__a21o_1 _13008_ (.A1(_05687_),
    .A2(_05695_),
    .B1(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__xor2_1 _13009_ (.A(_05666_),
    .B(_05697_),
    .X(_05698_));
 sky130_fd_sc_hd__clkinv_2 _13010_ (.A(_05671_),
    .Y(_05699_));
 sky130_fd_sc_hd__nor2_2 _13011_ (.A(_05433_),
    .B(_05606_),
    .Y(_05700_));
 sky130_fd_sc_hd__buf_2 _13012_ (.A(_05700_),
    .X(_05701_));
 sky130_fd_sc_hd__or2_1 _13013_ (.A(_05604_),
    .B(_05582_),
    .X(_05702_));
 sky130_fd_sc_hd__or3b_4 _13014_ (.A(_05591_),
    .B(_05702_),
    .C_N(_05566_),
    .X(_05703_));
 sky130_fd_sc_hd__a21o_1 _13015_ (.A1(_05566_),
    .A2(_05605_),
    .B1(_05583_),
    .X(_05704_));
 sky130_fd_sc_hd__a21o_1 _13016_ (.A1(_05703_),
    .A2(_05704_),
    .B1(_05629_),
    .X(_05705_));
 sky130_fd_sc_hd__nand2_1 _13017_ (.A(_05567_),
    .B(_05605_),
    .Y(_05706_));
 sky130_fd_sc_hd__a21bo_1 _13018_ (.A1(_05645_),
    .A2(_05567_),
    .B1_N(_05604_),
    .X(_05707_));
 sky130_fd_sc_hd__a21oi_1 _13019_ (.A1(_05706_),
    .A2(_05707_),
    .B1(_05625_),
    .Y(_05708_));
 sky130_fd_sc_hd__xnor2_1 _13020_ (.A(_05705_),
    .B(_05708_),
    .Y(_05709_));
 sky130_fd_sc_hd__nand2_1 _13021_ (.A(_05703_),
    .B(_05704_),
    .Y(_05710_));
 sky130_fd_sc_hd__and3_1 _13022_ (.A(_05612_),
    .B(_05710_),
    .C(_05708_),
    .X(_05711_));
 sky130_fd_sc_hd__a31o_1 _13023_ (.A1(_05699_),
    .A2(_05701_),
    .A3(_05709_),
    .B1(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__nand2_1 _13024_ (.A(_05612_),
    .B(_05700_),
    .Y(_05713_));
 sky130_fd_sc_hd__a21o_1 _13025_ (.A1(_05703_),
    .A2(_05704_),
    .B1(_05625_),
    .X(_05714_));
 sky130_fd_sc_hd__buf_2 _13026_ (.A(_05635_),
    .X(_05715_));
 sky130_fd_sc_hd__a21oi_1 _13027_ (.A1(_05706_),
    .A2(_05707_),
    .B1(_05715_),
    .Y(_05716_));
 sky130_fd_sc_hd__xnor2_1 _13028_ (.A(_05714_),
    .B(_05716_),
    .Y(_05717_));
 sky130_fd_sc_hd__xnor2_2 _13029_ (.A(_05713_),
    .B(_05717_),
    .Y(_05718_));
 sky130_fd_sc_hd__nand2_1 _13030_ (.A(_05712_),
    .B(_05718_),
    .Y(_05719_));
 sky130_fd_sc_hd__and2b_1 _13031_ (.A_N(_05691_),
    .B(_05694_),
    .X(_05720_));
 sky130_fd_sc_hd__a21o_1 _13032_ (.A1(_05688_),
    .A2(_05690_),
    .B1(_05720_),
    .X(_05721_));
 sky130_fd_sc_hd__clkbuf_2 _13033_ (.A(_05710_),
    .X(_05722_));
 sky130_fd_sc_hd__and3_1 _13034_ (.A(_05525_),
    .B(_05722_),
    .C(_05716_),
    .X(_05723_));
 sky130_fd_sc_hd__a31o_1 _13035_ (.A1(_05612_),
    .A2(_05701_),
    .A3(_05717_),
    .B1(_05723_),
    .X(_05724_));
 sky130_fd_sc_hd__nand2_1 _13036_ (.A(_05525_),
    .B(_05700_),
    .Y(_05725_));
 sky130_fd_sc_hd__and2_1 _13037_ (.A(_05706_),
    .B(_05707_),
    .X(_05726_));
 sky130_fd_sc_hd__and2_1 _13038_ (.A(_05703_),
    .B(_05704_),
    .X(_05727_));
 sky130_fd_sc_hd__clkbuf_2 _13039_ (.A(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__or2_1 _13040_ (.A(_05607_),
    .B(_05728_),
    .X(_05729_));
 sky130_fd_sc_hd__o22ai_1 _13041_ (.A1(_05715_),
    .A2(_05728_),
    .B1(_05726_),
    .B2(_05607_),
    .Y(_05730_));
 sky130_fd_sc_hd__o31a_1 _13042_ (.A1(_05715_),
    .A2(_05726_),
    .A3(_05729_),
    .B1(_05730_),
    .X(_05731_));
 sky130_fd_sc_hd__xnor2_1 _13043_ (.A(_05725_),
    .B(_05731_),
    .Y(_05732_));
 sky130_fd_sc_hd__xor2_1 _13044_ (.A(_05724_),
    .B(_05732_),
    .X(_05733_));
 sky130_fd_sc_hd__xnor2_1 _13045_ (.A(_05721_),
    .B(_05733_),
    .Y(_05734_));
 sky130_fd_sc_hd__xnor2_1 _13046_ (.A(_05719_),
    .B(_05734_),
    .Y(_05735_));
 sky130_fd_sc_hd__or2b_1 _13047_ (.A(_05666_),
    .B_N(_05697_),
    .X(_05736_));
 sky130_fd_sc_hd__o21ai_1 _13048_ (.A1(_05698_),
    .A2(_05735_),
    .B1(_05736_),
    .Y(_05737_));
 sky130_fd_sc_hd__nand2_4 _13049_ (.A(_05634_),
    .B(_05636_),
    .Y(_05738_));
 sky130_fd_sc_hd__and3_1 _13050_ (.A(_05401_),
    .B(_05738_),
    .C(_05652_),
    .X(_05739_));
 sky130_fd_sc_hd__clkbuf_4 _13051_ (.A(_05622_),
    .X(_05740_));
 sky130_fd_sc_hd__o22a_1 _13052_ (.A1(_05433_),
    .A2(_05740_),
    .B1(_05638_),
    .B2(_05624_),
    .X(_05741_));
 sky130_fd_sc_hd__or2_1 _13053_ (.A(_05739_),
    .B(_05741_),
    .X(_05742_));
 sky130_fd_sc_hd__nor2_1 _13054_ (.A(_05608_),
    .B(_05619_),
    .Y(_05743_));
 sky130_fd_sc_hd__a21bo_1 _13055_ (.A1(_05653_),
    .A2(_05655_),
    .B1_N(_05642_),
    .X(_05744_));
 sky130_fd_sc_hd__a21o_2 _13056_ (.A1(_05526_),
    .A2(_05546_),
    .B1(_05553_),
    .X(_05745_));
 sky130_fd_sc_hd__and2_1 _13057_ (.A(_05618_),
    .B(_05745_),
    .X(_05746_));
 sky130_fd_sc_hd__nor2_1 _13058_ (.A(_05621_),
    .B(_05746_),
    .Y(_05747_));
 sky130_fd_sc_hd__or4_4 _13059_ (.A(_05564_),
    .B(_05613_),
    .C(_05614_),
    .D(_05616_),
    .X(_05748_));
 sky130_fd_sc_hd__nand2_2 _13060_ (.A(_05567_),
    .B(_05748_),
    .Y(_05749_));
 sky130_fd_sc_hd__nor2_1 _13061_ (.A(_05608_),
    .B(_05749_),
    .Y(_05750_));
 sky130_fd_sc_hd__xor2_1 _13062_ (.A(_05747_),
    .B(_05750_),
    .X(_05751_));
 sky130_fd_sc_hd__nor2_1 _13063_ (.A(_05608_),
    .B(_05611_),
    .Y(_05752_));
 sky130_fd_sc_hd__xnor2_1 _13064_ (.A(_05751_),
    .B(_05752_),
    .Y(_05753_));
 sky130_fd_sc_hd__xnor2_1 _13065_ (.A(_05744_),
    .B(_05753_),
    .Y(_05754_));
 sky130_fd_sc_hd__xnor2_1 _13066_ (.A(_05743_),
    .B(_05754_),
    .Y(_05755_));
 sky130_fd_sc_hd__nor2_1 _13067_ (.A(_05742_),
    .B(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__and2_1 _13068_ (.A(_05742_),
    .B(_05755_),
    .X(_05757_));
 sky130_fd_sc_hd__or2_1 _13069_ (.A(_05756_),
    .B(_05757_),
    .X(_05758_));
 sky130_fd_sc_hd__or2b_1 _13070_ (.A(_05656_),
    .B_N(_05664_),
    .X(_05759_));
 sky130_fd_sc_hd__a21bo_1 _13071_ (.A1(_05650_),
    .A2(_05665_),
    .B1_N(_05759_),
    .X(_05760_));
 sky130_fd_sc_hd__xnor2_1 _13072_ (.A(_05758_),
    .B(_05760_),
    .Y(_05761_));
 sky130_fd_sc_hd__nand2_1 _13073_ (.A(_05724_),
    .B(_05732_),
    .Y(_05762_));
 sky130_fd_sc_hd__and2b_1 _13074_ (.A_N(_05648_),
    .B(_05644_),
    .X(_05763_));
 sky130_fd_sc_hd__and2b_1 _13075_ (.A_N(_05620_),
    .B(_05649_),
    .X(_05764_));
 sky130_fd_sc_hd__or2_1 _13076_ (.A(_05763_),
    .B(_05764_),
    .X(_05765_));
 sky130_fd_sc_hd__inv_2 _13077_ (.A(_05635_),
    .Y(_05766_));
 sky130_fd_sc_hd__buf_2 _13078_ (.A(_05726_),
    .X(_05767_));
 sky130_fd_sc_hd__nor2_1 _13079_ (.A(_05607_),
    .B(_05767_),
    .Y(_05768_));
 sky130_fd_sc_hd__and3_1 _13080_ (.A(_05766_),
    .B(_05722_),
    .C(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__and3_1 _13081_ (.A(_05525_),
    .B(_05701_),
    .C(_05731_),
    .X(_05770_));
 sky130_fd_sc_hd__nand2_1 _13082_ (.A(_05766_),
    .B(_05700_),
    .Y(_05771_));
 sky130_fd_sc_hd__nor2_1 _13083_ (.A(_05616_),
    .B(_05726_),
    .Y(_05772_));
 sky130_fd_sc_hd__xnor2_1 _13084_ (.A(_05729_),
    .B(_05772_),
    .Y(_05773_));
 sky130_fd_sc_hd__xnor2_1 _13085_ (.A(_05771_),
    .B(_05773_),
    .Y(_05774_));
 sky130_fd_sc_hd__o21ai_2 _13086_ (.A1(_05769_),
    .A2(_05770_),
    .B1(_05774_),
    .Y(_05775_));
 sky130_fd_sc_hd__or3_1 _13087_ (.A(_05769_),
    .B(_05770_),
    .C(_05774_),
    .X(_05776_));
 sky130_fd_sc_hd__and2_1 _13088_ (.A(_05775_),
    .B(_05776_),
    .X(_05777_));
 sky130_fd_sc_hd__xnor2_1 _13089_ (.A(_05765_),
    .B(_05777_),
    .Y(_05778_));
 sky130_fd_sc_hd__xor2_1 _13090_ (.A(_05762_),
    .B(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__xnor2_1 _13091_ (.A(_05761_),
    .B(_05779_),
    .Y(_05780_));
 sky130_fd_sc_hd__xnor2_1 _13092_ (.A(_05737_),
    .B(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__nand2_1 _13093_ (.A(_05721_),
    .B(_05733_),
    .Y(_05782_));
 sky130_fd_sc_hd__o21a_1 _13094_ (.A1(_05719_),
    .A2(_05734_),
    .B1(_05782_),
    .X(_05783_));
 sky130_fd_sc_hd__xor2_1 _13095_ (.A(_05781_),
    .B(_05783_),
    .X(_05784_));
 sky130_fd_sc_hd__a21oi_1 _13096_ (.A1(_05682_),
    .A2(_05683_),
    .B1(_05684_),
    .Y(_05785_));
 sky130_fd_sc_hd__nor2_1 _13097_ (.A(_05685_),
    .B(_05785_),
    .Y(_05786_));
 sky130_fd_sc_hd__a21oi_1 _13098_ (.A1(_05692_),
    .A2(_05641_),
    .B1(_05679_),
    .Y(_05787_));
 sky130_fd_sc_hd__and3_1 _13099_ (.A(_05692_),
    .B(_05640_),
    .C(_05679_),
    .X(_05788_));
 sky130_fd_sc_hd__nor2_1 _13100_ (.A(_05787_),
    .B(_05788_),
    .Y(_05789_));
 sky130_fd_sc_hd__nor2_1 _13101_ (.A(_05616_),
    .B(_05638_),
    .Y(_05790_));
 sky130_fd_sc_hd__xor2_1 _13102_ (.A(_05789_),
    .B(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__xor2_1 _13103_ (.A(_05674_),
    .B(_05675_),
    .X(_05792_));
 sky130_fd_sc_hd__buf_2 _13104_ (.A(_05672_),
    .X(_05793_));
 sky130_fd_sc_hd__nor3_1 _13105_ (.A(_05793_),
    .B(_05621_),
    .C(_05658_),
    .Y(_05794_));
 sky130_fd_sc_hd__or2_1 _13106_ (.A(_05608_),
    .B(_05660_),
    .X(_05795_));
 sky130_fd_sc_hd__or3_1 _13107_ (.A(_05627_),
    .B(_05604_),
    .C(_05657_),
    .X(_05796_));
 sky130_fd_sc_hd__xor2_1 _13108_ (.A(_05673_),
    .B(_05796_),
    .X(_05797_));
 sky130_fd_sc_hd__nor2_1 _13109_ (.A(_05795_),
    .B(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__or3_1 _13110_ (.A(_05792_),
    .B(_05794_),
    .C(_05798_),
    .X(_05799_));
 sky130_fd_sc_hd__o21a_1 _13111_ (.A1(_05794_),
    .A2(_05798_),
    .B1(_05792_),
    .X(_05800_));
 sky130_fd_sc_hd__a21o_1 _13112_ (.A1(_05791_),
    .A2(_05799_),
    .B1(_05800_),
    .X(_05801_));
 sky130_fd_sc_hd__xnor2_1 _13113_ (.A(_05786_),
    .B(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__nor2_1 _13114_ (.A(_05625_),
    .B(_05609_),
    .Y(_05803_));
 sky130_fd_sc_hd__a21o_1 _13115_ (.A1(_05618_),
    .A2(_05745_),
    .B1(_05537_),
    .X(_05804_));
 sky130_fd_sc_hd__and3_1 _13116_ (.A(_05766_),
    .B(_05567_),
    .C(_05748_),
    .X(_05805_));
 sky130_fd_sc_hd__xnor2_1 _13117_ (.A(_05804_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__or3_1 _13118_ (.A(_05715_),
    .B(_05804_),
    .C(_05749_),
    .X(_05807_));
 sky130_fd_sc_hd__a21bo_1 _13119_ (.A1(_05803_),
    .A2(_05806_),
    .B1_N(_05807_),
    .X(_05808_));
 sky130_fd_sc_hd__a21oi_1 _13120_ (.A1(_05789_),
    .A2(_05790_),
    .B1(_05788_),
    .Y(_05809_));
 sky130_fd_sc_hd__o22ai_1 _13121_ (.A1(_05611_),
    .A2(_05607_),
    .B1(_05715_),
    .B2(_05610_),
    .Y(_05810_));
 sky130_fd_sc_hd__and2_1 _13122_ (.A(_05693_),
    .B(_05810_),
    .X(_05811_));
 sky130_fd_sc_hd__xnor2_1 _13123_ (.A(_05809_),
    .B(_05811_),
    .Y(_05812_));
 sky130_fd_sc_hd__xnor2_1 _13124_ (.A(_05808_),
    .B(_05812_),
    .Y(_05813_));
 sky130_fd_sc_hd__nand2_1 _13125_ (.A(_05786_),
    .B(_05801_),
    .Y(_05814_));
 sky130_fd_sc_hd__o21a_1 _13126_ (.A1(_05802_),
    .A2(_05813_),
    .B1(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__xnor2_1 _13127_ (.A(_05687_),
    .B(_05695_),
    .Y(_05816_));
 sky130_fd_sc_hd__xor2_1 _13128_ (.A(_05815_),
    .B(_05816_),
    .X(_05817_));
 sky130_fd_sc_hd__nand2_2 _13129_ (.A(_05706_),
    .B(_05707_),
    .Y(_05818_));
 sky130_fd_sc_hd__nand2_1 _13130_ (.A(_05699_),
    .B(_05818_),
    .Y(_05819_));
 sky130_fd_sc_hd__nand2_1 _13131_ (.A(_05488_),
    .B(_05700_),
    .Y(_05820_));
 sky130_fd_sc_hd__o22a_1 _13132_ (.A1(_05671_),
    .A2(_05728_),
    .B1(_05726_),
    .B2(_05629_),
    .X(_05821_));
 sky130_fd_sc_hd__o22a_1 _13133_ (.A1(_05705_),
    .A2(_05819_),
    .B1(_05820_),
    .B2(_05821_),
    .X(_05822_));
 sky130_fd_sc_hd__nand2_1 _13134_ (.A(_05699_),
    .B(_05700_),
    .Y(_05823_));
 sky130_fd_sc_hd__xnor2_1 _13135_ (.A(_05823_),
    .B(_05709_),
    .Y(_05824_));
 sky130_fd_sc_hd__or2b_1 _13136_ (.A(_05822_),
    .B_N(_05824_),
    .X(_05825_));
 sky130_fd_sc_hd__and2b_1 _13137_ (.A_N(_05809_),
    .B(_05811_),
    .X(_05826_));
 sky130_fd_sc_hd__a21o_1 _13138_ (.A1(_05808_),
    .A2(_05812_),
    .B1(_05826_),
    .X(_05827_));
 sky130_fd_sc_hd__xor2_1 _13139_ (.A(_05712_),
    .B(_05718_),
    .X(_05828_));
 sky130_fd_sc_hd__xnor2_1 _13140_ (.A(_05827_),
    .B(_05828_),
    .Y(_05829_));
 sky130_fd_sc_hd__xor2_1 _13141_ (.A(_05825_),
    .B(_05829_),
    .X(_05830_));
 sky130_fd_sc_hd__nor2_1 _13142_ (.A(_05815_),
    .B(_05816_),
    .Y(_05831_));
 sky130_fd_sc_hd__a21o_1 _13143_ (.A1(_05817_),
    .A2(_05830_),
    .B1(_05831_),
    .X(_05832_));
 sky130_fd_sc_hd__xor2_1 _13144_ (.A(_05698_),
    .B(_05735_),
    .X(_05833_));
 sky130_fd_sc_hd__xnor2_1 _13145_ (.A(_05832_),
    .B(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__nand2_1 _13146_ (.A(_05827_),
    .B(_05828_),
    .Y(_05835_));
 sky130_fd_sc_hd__o21a_1 _13147_ (.A1(_05825_),
    .A2(_05829_),
    .B1(_05835_),
    .X(_05836_));
 sky130_fd_sc_hd__nand2_1 _13148_ (.A(_05832_),
    .B(_05833_),
    .Y(_05837_));
 sky130_fd_sc_hd__o21ai_1 _13149_ (.A1(_05834_),
    .A2(_05836_),
    .B1(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__nor2b_1 _13150_ (.A(_05784_),
    .B_N(_05838_),
    .Y(_05839_));
 sky130_fd_sc_hd__or2b_1 _13151_ (.A(_05780_),
    .B_N(_05737_),
    .X(_05840_));
 sky130_fd_sc_hd__or2b_1 _13152_ (.A(_05783_),
    .B_N(_05781_),
    .X(_05841_));
 sky130_fd_sc_hd__nand2_1 _13153_ (.A(_05840_),
    .B(_05841_),
    .Y(_05842_));
 sky130_fd_sc_hd__and2b_1 _13154_ (.A_N(_05758_),
    .B(_05760_),
    .X(_05843_));
 sky130_fd_sc_hd__and2_1 _13155_ (.A(_05761_),
    .B(_05779_),
    .X(_05844_));
 sky130_fd_sc_hd__nand2_1 _13156_ (.A(_05401_),
    .B(_05738_),
    .Y(_05845_));
 sky130_fd_sc_hd__a22o_1 _13157_ (.A1(_05747_),
    .A2(_05750_),
    .B1(_05751_),
    .B2(_05752_),
    .X(_05846_));
 sky130_fd_sc_hd__and2_1 _13158_ (.A(_05645_),
    .B(_05567_),
    .X(_05847_));
 sky130_fd_sc_hd__nor2_1 _13159_ (.A(_05624_),
    .B(_05749_),
    .Y(_05848_));
 sky130_fd_sc_hd__and2_1 _13160_ (.A(_05747_),
    .B(_05848_),
    .X(_05849_));
 sky130_fd_sc_hd__o22a_1 _13161_ (.A1(_05624_),
    .A2(_05746_),
    .B1(_05749_),
    .B2(_05621_),
    .X(_05850_));
 sky130_fd_sc_hd__or2_1 _13162_ (.A(_05849_),
    .B(_05850_),
    .X(_05851_));
 sky130_fd_sc_hd__xnor2_1 _13163_ (.A(_05847_),
    .B(_05851_),
    .Y(_05852_));
 sky130_fd_sc_hd__xnor2_1 _13164_ (.A(_05739_),
    .B(_05852_),
    .Y(_05853_));
 sky130_fd_sc_hd__xnor2_1 _13165_ (.A(_05846_),
    .B(_05853_),
    .Y(_05854_));
 sky130_fd_sc_hd__xnor2_1 _13166_ (.A(_05845_),
    .B(_05854_),
    .Y(_05855_));
 sky130_fd_sc_hd__xnor2_1 _13167_ (.A(_05756_),
    .B(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__or2b_1 _13168_ (.A(_05753_),
    .B_N(_05744_),
    .X(_05857_));
 sky130_fd_sc_hd__a21bo_1 _13169_ (.A1(_05743_),
    .A2(_05754_),
    .B1_N(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__and3_1 _13170_ (.A(_05553_),
    .B(_05722_),
    .C(_05768_),
    .X(_05859_));
 sky130_fd_sc_hd__and3_1 _13171_ (.A(_05766_),
    .B(_05701_),
    .C(_05773_),
    .X(_05860_));
 sky130_fd_sc_hd__nand2_4 _13172_ (.A(_05401_),
    .B(_05703_),
    .Y(_05861_));
 sky130_fd_sc_hd__or2_1 _13173_ (.A(_05607_),
    .B(_05861_),
    .X(_05862_));
 sky130_fd_sc_hd__o22a_1 _13174_ (.A1(_05616_),
    .A2(_05728_),
    .B1(_05726_),
    .B2(_05611_),
    .X(_05863_));
 sky130_fd_sc_hd__a31oi_1 _13175_ (.A1(_05692_),
    .A2(_05710_),
    .A3(_05772_),
    .B1(_05863_),
    .Y(_05864_));
 sky130_fd_sc_hd__xnor2_1 _13176_ (.A(_05862_),
    .B(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__o21ai_1 _13177_ (.A1(_05859_),
    .A2(_05860_),
    .B1(_05865_),
    .Y(_05866_));
 sky130_fd_sc_hd__or3_1 _13178_ (.A(_05859_),
    .B(_05860_),
    .C(_05865_),
    .X(_05867_));
 sky130_fd_sc_hd__and2_1 _13179_ (.A(_05866_),
    .B(_05867_),
    .X(_05868_));
 sky130_fd_sc_hd__xnor2_1 _13180_ (.A(_05858_),
    .B(_05868_),
    .Y(_05869_));
 sky130_fd_sc_hd__xor2_1 _13181_ (.A(_05775_),
    .B(_05869_),
    .X(_05870_));
 sky130_fd_sc_hd__xnor2_1 _13182_ (.A(_05856_),
    .B(_05870_),
    .Y(_05871_));
 sky130_fd_sc_hd__o21ai_1 _13183_ (.A1(_05843_),
    .A2(_05844_),
    .B1(_05871_),
    .Y(_05872_));
 sky130_fd_sc_hd__or3_1 _13184_ (.A(_05843_),
    .B(_05844_),
    .C(_05871_),
    .X(_05873_));
 sky130_fd_sc_hd__and2_1 _13185_ (.A(_05872_),
    .B(_05873_),
    .X(_05874_));
 sky130_fd_sc_hd__nor2_1 _13186_ (.A(_05762_),
    .B(_05778_),
    .Y(_05875_));
 sky130_fd_sc_hd__a21oi_1 _13187_ (.A1(_05765_),
    .A2(_05777_),
    .B1(_05875_),
    .Y(_05876_));
 sky130_fd_sc_hd__xor2_1 _13188_ (.A(_05874_),
    .B(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__xnor2_1 _13189_ (.A(_05842_),
    .B(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__xor2_1 _13190_ (.A(_05839_),
    .B(_05878_),
    .X(_05879_));
 sky130_fd_sc_hd__and2b_1 _13191_ (.A_N(_05838_),
    .B(_05784_),
    .X(_05880_));
 sky130_fd_sc_hd__nor2_1 _13192_ (.A(_05839_),
    .B(_05880_),
    .Y(_05881_));
 sky130_fd_sc_hd__o21bai_1 _13193_ (.A1(_05705_),
    .A2(_05819_),
    .B1_N(_05821_),
    .Y(_05882_));
 sky130_fd_sc_hd__xnor2_2 _13194_ (.A(_05820_),
    .B(_05882_),
    .Y(_05883_));
 sky130_fd_sc_hd__or3_2 _13195_ (.A(_05793_),
    .B(_05728_),
    .C(_05819_),
    .X(_05884_));
 sky130_fd_sc_hd__xnor2_1 _13196_ (.A(_05822_),
    .B(_05824_),
    .Y(_05885_));
 sky130_fd_sc_hd__a21oi_1 _13197_ (.A1(_05626_),
    .A2(_05630_),
    .B1(_05616_),
    .Y(_05886_));
 sky130_fd_sc_hd__a22o_1 _13198_ (.A1(_05553_),
    .A2(_05640_),
    .B1(_05651_),
    .B2(_05692_),
    .X(_05887_));
 sky130_fd_sc_hd__or3b_1 _13199_ (.A(_05564_),
    .B(_05622_),
    .C_N(_05886_),
    .X(_05888_));
 sky130_fd_sc_hd__and3_1 _13200_ (.A(_05615_),
    .B(_05887_),
    .C(_05888_),
    .X(_05889_));
 sky130_fd_sc_hd__a31o_1 _13201_ (.A1(_05692_),
    .A2(_05641_),
    .A3(_05886_),
    .B1(_05889_),
    .X(_05890_));
 sky130_fd_sc_hd__xor2_1 _13202_ (.A(_05803_),
    .B(_05806_),
    .X(_05891_));
 sky130_fd_sc_hd__xnor2_1 _13203_ (.A(_05890_),
    .B(_05891_),
    .Y(_05892_));
 sky130_fd_sc_hd__a21o_1 _13204_ (.A1(_05618_),
    .A2(_05745_),
    .B1(_05625_),
    .X(_05893_));
 sky130_fd_sc_hd__or2_1 _13205_ (.A(_05629_),
    .B(_05609_),
    .X(_05894_));
 sky130_fd_sc_hd__a21o_1 _13206_ (.A1(_05618_),
    .A2(_05745_),
    .B1(_05635_),
    .X(_05895_));
 sky130_fd_sc_hd__and3_1 _13207_ (.A(_05525_),
    .B(_05567_),
    .C(_05748_),
    .X(_05896_));
 sky130_fd_sc_hd__xnor2_1 _13208_ (.A(_05895_),
    .B(_05896_),
    .Y(_05897_));
 sky130_fd_sc_hd__or2b_1 _13209_ (.A(_05894_),
    .B_N(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__o31a_1 _13210_ (.A1(_05715_),
    .A2(_05749_),
    .A3(_05893_),
    .B1(_05898_),
    .X(_05899_));
 sky130_fd_sc_hd__nand2_1 _13211_ (.A(_05890_),
    .B(_05891_),
    .Y(_05900_));
 sky130_fd_sc_hd__o21a_1 _13212_ (.A1(_05892_),
    .A2(_05899_),
    .B1(_05900_),
    .X(_05901_));
 sky130_fd_sc_hd__xor2_1 _13213_ (.A(_05885_),
    .B(_05901_),
    .X(_05902_));
 sky130_fd_sc_hd__or2b_1 _13214_ (.A(_05901_),
    .B_N(_05885_),
    .X(_05903_));
 sky130_fd_sc_hd__o31a_1 _13215_ (.A1(_05883_),
    .A2(_05884_),
    .A3(_05902_),
    .B1(_05903_),
    .X(_05904_));
 sky130_fd_sc_hd__xnor2_1 _13216_ (.A(_05817_),
    .B(_05830_),
    .Y(_05905_));
 sky130_fd_sc_hd__xnor2_1 _13217_ (.A(_05802_),
    .B(_05813_),
    .Y(_05906_));
 sky130_fd_sc_hd__xor2_1 _13218_ (.A(_05892_),
    .B(_05899_),
    .X(_05907_));
 sky130_fd_sc_hd__and2b_1 _13219_ (.A_N(_05800_),
    .B(_05799_),
    .X(_05908_));
 sky130_fd_sc_hd__xor2_1 _13220_ (.A(_05791_),
    .B(_05908_),
    .X(_05909_));
 sky130_fd_sc_hd__xnor2_1 _13221_ (.A(_05795_),
    .B(_05797_),
    .Y(_05910_));
 sky130_fd_sc_hd__or2_1 _13222_ (.A(_05591_),
    .B(_05672_),
    .X(_05911_));
 sky130_fd_sc_hd__nor2_1 _13223_ (.A(_05611_),
    .B(_05660_),
    .Y(_05912_));
 sky130_fd_sc_hd__nor2_1 _13224_ (.A(_05672_),
    .B(_05604_),
    .Y(_05913_));
 sky130_fd_sc_hd__or3_1 _13225_ (.A(_05591_),
    .B(_05627_),
    .C(_05657_),
    .X(_05914_));
 sky130_fd_sc_hd__xnor2_1 _13226_ (.A(_05913_),
    .B(_05914_),
    .Y(_05915_));
 sky130_fd_sc_hd__a2bb2o_1 _13227_ (.A1_N(_05796_),
    .A2_N(_05911_),
    .B1(_05912_),
    .B2(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__and2b_1 _13228_ (.A_N(_05910_),
    .B(_05916_),
    .X(_05917_));
 sky130_fd_sc_hd__xor2_1 _13229_ (.A(_05910_),
    .B(_05916_),
    .X(_05918_));
 sky130_fd_sc_hd__a21oi_1 _13230_ (.A1(_05887_),
    .A2(_05888_),
    .B1(_05615_),
    .Y(_05919_));
 sky130_fd_sc_hd__nor3_1 _13231_ (.A(_05918_),
    .B(_05889_),
    .C(_05919_),
    .Y(_05920_));
 sky130_fd_sc_hd__nor2_1 _13232_ (.A(_05917_),
    .B(_05920_),
    .Y(_05921_));
 sky130_fd_sc_hd__xnor2_1 _13233_ (.A(_05909_),
    .B(_05921_),
    .Y(_05922_));
 sky130_fd_sc_hd__and2b_1 _13234_ (.A_N(_05921_),
    .B(_05909_),
    .X(_05923_));
 sky130_fd_sc_hd__a21oi_1 _13235_ (.A1(_05907_),
    .A2(_05922_),
    .B1(_05923_),
    .Y(_05924_));
 sky130_fd_sc_hd__nand2_1 _13236_ (.A(_05906_),
    .B(_05924_),
    .Y(_05925_));
 sky130_fd_sc_hd__nor2_1 _13237_ (.A(_05883_),
    .B(_05884_),
    .Y(_05926_));
 sky130_fd_sc_hd__xnor2_1 _13238_ (.A(_05926_),
    .B(_05902_),
    .Y(_05927_));
 sky130_fd_sc_hd__nor2_1 _13239_ (.A(_05906_),
    .B(_05924_),
    .Y(_05928_));
 sky130_fd_sc_hd__a21oi_1 _13240_ (.A1(_05925_),
    .A2(_05927_),
    .B1(_05928_),
    .Y(_05929_));
 sky130_fd_sc_hd__xnor2_1 _13241_ (.A(_05905_),
    .B(_05929_),
    .Y(_05930_));
 sky130_fd_sc_hd__or2_1 _13242_ (.A(_05905_),
    .B(_05929_),
    .X(_05931_));
 sky130_fd_sc_hd__o21a_1 _13243_ (.A1(_05904_),
    .A2(_05930_),
    .B1(_05931_),
    .X(_05932_));
 sky130_fd_sc_hd__xor2_1 _13244_ (.A(_05834_),
    .B(_05836_),
    .X(_05933_));
 sky130_fd_sc_hd__and2b_1 _13245_ (.A_N(_05932_),
    .B(_05933_),
    .X(_05934_));
 sky130_fd_sc_hd__and2_1 _13246_ (.A(_05881_),
    .B(_05934_),
    .X(_05935_));
 sky130_fd_sc_hd__xor2_1 _13247_ (.A(_05879_),
    .B(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__xnor2_1 _13248_ (.A(_05904_),
    .B(_05930_),
    .Y(_05937_));
 sky130_fd_sc_hd__xnor2_1 _13249_ (.A(_05883_),
    .B(_05884_),
    .Y(_05938_));
 sky130_fd_sc_hd__xnor2_1 _13250_ (.A(_05894_),
    .B(_05897_),
    .Y(_05939_));
 sky130_fd_sc_hd__xnor2_1 _13251_ (.A(_05615_),
    .B(_05939_),
    .Y(_05940_));
 sky130_fd_sc_hd__a21oi_1 _13252_ (.A1(_05618_),
    .A2(_05745_),
    .B1(_05629_),
    .Y(_05941_));
 sky130_fd_sc_hd__nor2_1 _13253_ (.A(_05671_),
    .B(_05610_),
    .Y(_05942_));
 sky130_fd_sc_hd__and3_1 _13254_ (.A(_05612_),
    .B(_05567_),
    .C(_05748_),
    .X(_05943_));
 sky130_fd_sc_hd__xnor2_1 _13255_ (.A(_05893_),
    .B(_05943_),
    .Y(_05944_));
 sky130_fd_sc_hd__a22o_1 _13256_ (.A1(_05896_),
    .A2(_05941_),
    .B1(_05942_),
    .B2(_05944_),
    .X(_05945_));
 sky130_fd_sc_hd__or2b_1 _13257_ (.A(_05940_),
    .B_N(_05945_),
    .X(_05946_));
 sky130_fd_sc_hd__a21bo_1 _13258_ (.A1(_05615_),
    .A2(_05939_),
    .B1_N(_05946_),
    .X(_05947_));
 sky130_fd_sc_hd__and2b_1 _13259_ (.A_N(_05938_),
    .B(_05947_),
    .X(_05948_));
 sky130_fd_sc_hd__xnor2_1 _13260_ (.A(_05906_),
    .B(_05924_),
    .Y(_05949_));
 sky130_fd_sc_hd__xnor2_1 _13261_ (.A(_05949_),
    .B(_05927_),
    .Y(_05950_));
 sky130_fd_sc_hd__xnor2_1 _13262_ (.A(_05947_),
    .B(_05938_),
    .Y(_05951_));
 sky130_fd_sc_hd__xor2_1 _13263_ (.A(_05907_),
    .B(_05922_),
    .X(_05952_));
 sky130_fd_sc_hd__xnor2_1 _13264_ (.A(_05940_),
    .B(_05945_),
    .Y(_05953_));
 sky130_fd_sc_hd__o21a_1 _13265_ (.A1(_05889_),
    .A2(_05919_),
    .B1(_05918_),
    .X(_05954_));
 sky130_fd_sc_hd__nor2_1 _13266_ (.A(_05920_),
    .B(_05954_),
    .Y(_05955_));
 sky130_fd_sc_hd__xnor2_1 _13267_ (.A(_05912_),
    .B(_05915_),
    .Y(_05956_));
 sky130_fd_sc_hd__or2_1 _13268_ (.A(_05564_),
    .B(_05672_),
    .X(_05957_));
 sky130_fd_sc_hd__or2_1 _13269_ (.A(_05616_),
    .B(_05659_),
    .X(_05958_));
 sky130_fd_sc_hd__or2_4 _13270_ (.A(_05627_),
    .B(_05657_),
    .X(_05959_));
 sky130_fd_sc_hd__o21a_1 _13271_ (.A1(_05611_),
    .A2(_05959_),
    .B1(_05911_),
    .X(_05960_));
 sky130_fd_sc_hd__o22a_1 _13272_ (.A1(_05914_),
    .A2(_05957_),
    .B1(_05958_),
    .B2(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__xor2_1 _13273_ (.A(_05956_),
    .B(_05961_),
    .X(_05962_));
 sky130_fd_sc_hd__or3_1 _13274_ (.A(_05537_),
    .B(_05622_),
    .C(_05886_),
    .X(_05963_));
 sky130_fd_sc_hd__o21ai_1 _13275_ (.A1(_05537_),
    .A2(_05622_),
    .B1(_05886_),
    .Y(_05964_));
 sky130_fd_sc_hd__a211o_1 _13276_ (.A1(_05963_),
    .A2(_05964_),
    .B1(_05635_),
    .C1(_05638_),
    .X(_05965_));
 sky130_fd_sc_hd__o211ai_1 _13277_ (.A1(_05715_),
    .A2(_05638_),
    .B1(_05963_),
    .C1(_05964_),
    .Y(_05966_));
 sky130_fd_sc_hd__and3_1 _13278_ (.A(_05962_),
    .B(_05965_),
    .C(_05966_),
    .X(_05967_));
 sky130_fd_sc_hd__o21ba_1 _13279_ (.A1(_05956_),
    .A2(_05961_),
    .B1_N(_05967_),
    .X(_05968_));
 sky130_fd_sc_hd__xnor2_1 _13280_ (.A(_05955_),
    .B(_05968_),
    .Y(_05969_));
 sky130_fd_sc_hd__and2b_1 _13281_ (.A_N(_05968_),
    .B(_05955_),
    .X(_05970_));
 sky130_fd_sc_hd__a21oi_1 _13282_ (.A1(_05953_),
    .A2(_05969_),
    .B1(_05970_),
    .Y(_05971_));
 sky130_fd_sc_hd__xnor2_1 _13283_ (.A(_05952_),
    .B(_05971_),
    .Y(_05972_));
 sky130_fd_sc_hd__and2b_1 _13284_ (.A_N(_05971_),
    .B(_05952_),
    .X(_05973_));
 sky130_fd_sc_hd__a21oi_1 _13285_ (.A1(_05951_),
    .A2(_05972_),
    .B1(_05973_),
    .Y(_05974_));
 sky130_fd_sc_hd__xnor2_1 _13286_ (.A(_05950_),
    .B(_05974_),
    .Y(_05975_));
 sky130_fd_sc_hd__or2b_1 _13287_ (.A(_05974_),
    .B_N(_05950_),
    .X(_05976_));
 sky130_fd_sc_hd__a21boi_1 _13288_ (.A1(_05948_),
    .A2(_05975_),
    .B1_N(_05976_),
    .Y(_05977_));
 sky130_fd_sc_hd__nor2_1 _13289_ (.A(_05937_),
    .B(_05977_),
    .Y(_05978_));
 sky130_fd_sc_hd__xnor2_1 _13290_ (.A(_05933_),
    .B(_05932_),
    .Y(_05979_));
 sky130_fd_sc_hd__and2_1 _13291_ (.A(_05978_),
    .B(_05979_),
    .X(_05980_));
 sky130_fd_sc_hd__xnor2_2 _13292_ (.A(_05948_),
    .B(_05975_),
    .Y(_05981_));
 sky130_fd_sc_hd__xnor2_1 _13293_ (.A(_05942_),
    .B(_05944_),
    .Y(_05982_));
 sky130_fd_sc_hd__nor2_1 _13294_ (.A(_05634_),
    .B(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__xnor2_1 _13295_ (.A(_05615_),
    .B(_05982_),
    .Y(_05984_));
 sky130_fd_sc_hd__and3_1 _13296_ (.A(_05699_),
    .B(_05567_),
    .C(_05748_),
    .X(_05985_));
 sky130_fd_sc_hd__nor2_1 _13297_ (.A(_05793_),
    .B(_05610_),
    .Y(_05986_));
 sky130_fd_sc_hd__xor2_1 _13298_ (.A(_05941_),
    .B(_05985_),
    .X(_05987_));
 sky130_fd_sc_hd__a22o_1 _13299_ (.A1(_05941_),
    .A2(_05985_),
    .B1(_05986_),
    .B2(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__and2_1 _13300_ (.A(_05984_),
    .B(_05988_),
    .X(_05989_));
 sky130_fd_sc_hd__o21ai_1 _13301_ (.A1(_05793_),
    .A2(_05728_),
    .B1(_05819_),
    .Y(_05990_));
 sky130_fd_sc_hd__and2_1 _13302_ (.A(_05884_),
    .B(_05990_),
    .X(_05991_));
 sky130_fd_sc_hd__o21a_1 _13303_ (.A1(_05983_),
    .A2(_05989_),
    .B1(_05991_),
    .X(_05992_));
 sky130_fd_sc_hd__xnor2_1 _13304_ (.A(_05951_),
    .B(_05972_),
    .Y(_05993_));
 sky130_fd_sc_hd__nor3_1 _13305_ (.A(_05983_),
    .B(_05989_),
    .C(_05991_),
    .Y(_05994_));
 sky130_fd_sc_hd__nor2_1 _13306_ (.A(_05992_),
    .B(_05994_),
    .Y(_05995_));
 sky130_fd_sc_hd__xnor2_1 _13307_ (.A(_05953_),
    .B(_05969_),
    .Y(_05996_));
 sky130_fd_sc_hd__xor2_1 _13308_ (.A(_05984_),
    .B(_05988_),
    .X(_05997_));
 sky130_fd_sc_hd__a21oi_1 _13309_ (.A1(_05965_),
    .A2(_05966_),
    .B1(_05962_),
    .Y(_05998_));
 sky130_fd_sc_hd__or2_1 _13310_ (.A(_05967_),
    .B(_05998_),
    .X(_05999_));
 sky130_fd_sc_hd__o21ba_1 _13311_ (.A1(_05914_),
    .A2(_05957_),
    .B1_N(_05960_),
    .X(_06000_));
 sky130_fd_sc_hd__xor2_1 _13312_ (.A(_05958_),
    .B(_06000_),
    .X(_06001_));
 sky130_fd_sc_hd__or3_2 _13313_ (.A(_05627_),
    .B(_05616_),
    .C(_05657_),
    .X(_06002_));
 sky130_fd_sc_hd__or2_1 _13314_ (.A(_05607_),
    .B(_05660_),
    .X(_06003_));
 sky130_fd_sc_hd__xnor2_1 _13315_ (.A(_05957_),
    .B(_06002_),
    .Y(_06004_));
 sky130_fd_sc_hd__o22ai_1 _13316_ (.A1(_05957_),
    .A2(_06002_),
    .B1(_06003_),
    .B2(_06004_),
    .Y(_06005_));
 sky130_fd_sc_hd__xor2_1 _13317_ (.A(_06001_),
    .B(_06005_),
    .X(_06006_));
 sky130_fd_sc_hd__nand2_1 _13318_ (.A(_05489_),
    .B(_05612_),
    .Y(_06007_));
 sky130_fd_sc_hd__or2_1 _13319_ (.A(_06007_),
    .B(_05635_),
    .X(_06008_));
 sky130_fd_sc_hd__nand2_1 _13320_ (.A(_05625_),
    .B(_06008_),
    .Y(_06009_));
 sky130_fd_sc_hd__or2_1 _13321_ (.A(_05607_),
    .B(_06007_),
    .X(_06010_));
 sky130_fd_sc_hd__xor2_1 _13322_ (.A(_06009_),
    .B(_06010_),
    .X(_06011_));
 sky130_fd_sc_hd__or2b_1 _13323_ (.A(_06001_),
    .B_N(_06005_),
    .X(_06012_));
 sky130_fd_sc_hd__o21a_1 _13324_ (.A1(_06006_),
    .A2(_06011_),
    .B1(_06012_),
    .X(_06013_));
 sky130_fd_sc_hd__xor2_1 _13325_ (.A(_05999_),
    .B(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__nor2_1 _13326_ (.A(_05999_),
    .B(_06013_),
    .Y(_06015_));
 sky130_fd_sc_hd__a21o_1 _13327_ (.A1(_05997_),
    .A2(_06014_),
    .B1(_06015_),
    .X(_06016_));
 sky130_fd_sc_hd__xnor2_1 _13328_ (.A(_05996_),
    .B(_06016_),
    .Y(_06017_));
 sky130_fd_sc_hd__or2b_1 _13329_ (.A(_05996_),
    .B_N(_06016_),
    .X(_06018_));
 sky130_fd_sc_hd__a21boi_1 _13330_ (.A1(_05995_),
    .A2(_06017_),
    .B1_N(_06018_),
    .Y(_06019_));
 sky130_fd_sc_hd__xor2_1 _13331_ (.A(_05993_),
    .B(_06019_),
    .X(_06020_));
 sky130_fd_sc_hd__nor2_1 _13332_ (.A(_05993_),
    .B(_06019_),
    .Y(_06021_));
 sky130_fd_sc_hd__a21oi_2 _13333_ (.A1(_05992_),
    .A2(_06020_),
    .B1(_06021_),
    .Y(_06022_));
 sky130_fd_sc_hd__nor2_1 _13334_ (.A(_05981_),
    .B(_06022_),
    .Y(_06023_));
 sky130_fd_sc_hd__xor2_1 _13335_ (.A(_05937_),
    .B(_05977_),
    .X(_06024_));
 sky130_fd_sc_hd__and2_1 _13336_ (.A(_06023_),
    .B(_06024_),
    .X(_06025_));
 sky130_fd_sc_hd__xor2_1 _13337_ (.A(_05981_),
    .B(_06022_),
    .X(_06026_));
 sky130_fd_sc_hd__xnor2_1 _13338_ (.A(_05995_),
    .B(_06017_),
    .Y(_06027_));
 sky130_fd_sc_hd__clkbuf_4 _13339_ (.A(_05488_),
    .X(_06028_));
 sky130_fd_sc_hd__nand2_1 _13340_ (.A(_06028_),
    .B(_05818_),
    .Y(_06029_));
 sky130_fd_sc_hd__xor2_1 _13341_ (.A(_05986_),
    .B(_05987_),
    .X(_06030_));
 sky130_fd_sc_hd__a21oi_1 _13342_ (.A1(_05626_),
    .A2(_06010_),
    .B1(_05715_),
    .Y(_06031_));
 sky130_fd_sc_hd__nor2_1 _13343_ (.A(_05671_),
    .B(_05746_),
    .Y(_06032_));
 sky130_fd_sc_hd__xor2_1 _13344_ (.A(_06030_),
    .B(_06031_),
    .X(_06033_));
 sky130_fd_sc_hd__nor2_1 _13345_ (.A(_05793_),
    .B(_05749_),
    .Y(_06034_));
 sky130_fd_sc_hd__and3_1 _13346_ (.A(_06032_),
    .B(_06033_),
    .C(_06034_),
    .X(_06035_));
 sky130_fd_sc_hd__a21oi_1 _13347_ (.A1(_06030_),
    .A2(_06031_),
    .B1(_06035_),
    .Y(_06036_));
 sky130_fd_sc_hd__xor2_1 _13348_ (.A(_06029_),
    .B(_06036_),
    .X(_06037_));
 sky130_fd_sc_hd__xor2_1 _13349_ (.A(_05997_),
    .B(_06014_),
    .X(_06038_));
 sky130_fd_sc_hd__nand2_1 _13350_ (.A(_06032_),
    .B(_06034_),
    .Y(_06039_));
 sky130_fd_sc_hd__xor2_1 _13351_ (.A(_06033_),
    .B(_06039_),
    .X(_06040_));
 sky130_fd_sc_hd__xor2_1 _13352_ (.A(_06006_),
    .B(_06011_),
    .X(_06041_));
 sky130_fd_sc_hd__or2_1 _13353_ (.A(_05537_),
    .B(_05793_),
    .X(_06042_));
 sky130_fd_sc_hd__or2_1 _13354_ (.A(_05635_),
    .B(_05660_),
    .X(_06043_));
 sky130_fd_sc_hd__or2_1 _13355_ (.A(_05793_),
    .B(_05616_),
    .X(_06044_));
 sky130_fd_sc_hd__or3_1 _13356_ (.A(_05537_),
    .B(_05627_),
    .C(_05657_),
    .X(_06045_));
 sky130_fd_sc_hd__xnor2_1 _13357_ (.A(_06044_),
    .B(_06045_),
    .Y(_06046_));
 sky130_fd_sc_hd__o22ai_2 _13358_ (.A1(_06002_),
    .A2(_06042_),
    .B1(_06043_),
    .B2(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__xnor2_1 _13359_ (.A(_06003_),
    .B(_06004_),
    .Y(_06048_));
 sky130_fd_sc_hd__or2b_1 _13360_ (.A(_06047_),
    .B_N(_06048_),
    .X(_06049_));
 sky130_fd_sc_hd__a21oi_1 _13361_ (.A1(_05634_),
    .A2(_05636_),
    .B1(_05629_),
    .Y(_06050_));
 sky130_fd_sc_hd__mux2_1 _13362_ (.A0(_05607_),
    .A1(_06050_),
    .S(_06008_),
    .X(_06051_));
 sky130_fd_sc_hd__and2b_1 _13363_ (.A_N(_06048_),
    .B(_06047_),
    .X(_06052_));
 sky130_fd_sc_hd__a21oi_1 _13364_ (.A1(_06049_),
    .A2(_06051_),
    .B1(_06052_),
    .Y(_06053_));
 sky130_fd_sc_hd__xor2_1 _13365_ (.A(_06041_),
    .B(_06053_),
    .X(_06054_));
 sky130_fd_sc_hd__or2b_1 _13366_ (.A(_06053_),
    .B_N(_06041_),
    .X(_06055_));
 sky130_fd_sc_hd__o21a_1 _13367_ (.A1(_06040_),
    .A2(_06054_),
    .B1(_06055_),
    .X(_06056_));
 sky130_fd_sc_hd__xnor2_1 _13368_ (.A(_06038_),
    .B(_06056_),
    .Y(_06057_));
 sky130_fd_sc_hd__and2b_1 _13369_ (.A_N(_06056_),
    .B(_06038_),
    .X(_06058_));
 sky130_fd_sc_hd__a21oi_1 _13370_ (.A1(_06037_),
    .A2(_06057_),
    .B1(_06058_),
    .Y(_06059_));
 sky130_fd_sc_hd__or2_1 _13371_ (.A(_06027_),
    .B(_06059_),
    .X(_06060_));
 sky130_fd_sc_hd__or2_1 _13372_ (.A(_06029_),
    .B(_06036_),
    .X(_06061_));
 sky130_fd_sc_hd__xor2_1 _13373_ (.A(_06027_),
    .B(_06059_),
    .X(_06062_));
 sky130_fd_sc_hd__or2b_1 _13374_ (.A(_06061_),
    .B_N(_06062_),
    .X(_06063_));
 sky130_fd_sc_hd__xnor2_1 _13375_ (.A(_05992_),
    .B(_06020_),
    .Y(_06064_));
 sky130_fd_sc_hd__a21oi_1 _13376_ (.A1(_06060_),
    .A2(_06063_),
    .B1(_06064_),
    .Y(_06065_));
 sky130_fd_sc_hd__xor2_1 _13377_ (.A(_06061_),
    .B(_06062_),
    .X(_06066_));
 sky130_fd_sc_hd__and3_1 _13378_ (.A(_06064_),
    .B(_06060_),
    .C(_06063_),
    .X(_06067_));
 sky130_fd_sc_hd__xnor2_1 _13379_ (.A(_06040_),
    .B(_06054_),
    .Y(_06068_));
 sky130_fd_sc_hd__xor2_1 _13380_ (.A(_06048_),
    .B(_06047_),
    .X(_06069_));
 sky130_fd_sc_hd__xnor2_1 _13381_ (.A(_06069_),
    .B(_06051_),
    .Y(_06070_));
 sky130_fd_sc_hd__or3_1 _13382_ (.A(_05629_),
    .B(_05715_),
    .C(_05626_),
    .X(_06071_));
 sky130_fd_sc_hd__o21ai_1 _13383_ (.A1(_05629_),
    .A2(_05622_),
    .B1(_05626_),
    .Y(_06072_));
 sky130_fd_sc_hd__nand4_2 _13384_ (.A(_05699_),
    .B(_05738_),
    .C(_06071_),
    .D(_06072_),
    .Y(_06073_));
 sky130_fd_sc_hd__a22o_1 _13385_ (.A1(_05699_),
    .A2(_05738_),
    .B1(_06071_),
    .B2(_06072_),
    .X(_06074_));
 sky130_fd_sc_hd__xnor2_1 _13386_ (.A(_06043_),
    .B(_06046_),
    .Y(_06075_));
 sky130_fd_sc_hd__or3_1 _13387_ (.A(_05627_),
    .B(_05635_),
    .C(_05657_),
    .X(_06076_));
 sky130_fd_sc_hd__or2_1 _13388_ (.A(_05625_),
    .B(_05660_),
    .X(_06077_));
 sky130_fd_sc_hd__xnor2_1 _13389_ (.A(_06042_),
    .B(_06076_),
    .Y(_06078_));
 sky130_fd_sc_hd__o22ai_2 _13390_ (.A1(_06042_),
    .A2(_06076_),
    .B1(_06077_),
    .B2(_06078_),
    .Y(_06079_));
 sky130_fd_sc_hd__xnor2_1 _13391_ (.A(_06075_),
    .B(_06079_),
    .Y(_06080_));
 sky130_fd_sc_hd__and2b_1 _13392_ (.A_N(_06075_),
    .B(_06079_),
    .X(_06081_));
 sky130_fd_sc_hd__a31o_1 _13393_ (.A1(_06073_),
    .A2(_06074_),
    .A3(_06080_),
    .B1(_06081_),
    .X(_06082_));
 sky130_fd_sc_hd__nand2_1 _13394_ (.A(_06071_),
    .B(_06073_),
    .Y(_06083_));
 sky130_fd_sc_hd__xnor2_1 _13395_ (.A(_06032_),
    .B(_06034_),
    .Y(_06084_));
 sky130_fd_sc_hd__xnor2_1 _13396_ (.A(_06083_),
    .B(_06084_),
    .Y(_06085_));
 sky130_fd_sc_hd__xor2_1 _13397_ (.A(_06070_),
    .B(_06082_),
    .X(_06086_));
 sky130_fd_sc_hd__nand2_1 _13398_ (.A(_06085_),
    .B(_06086_),
    .Y(_06087_));
 sky130_fd_sc_hd__a21bo_1 _13399_ (.A1(_06070_),
    .A2(_06082_),
    .B1_N(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__or2b_1 _13400_ (.A(_06068_),
    .B_N(_06088_),
    .X(_06089_));
 sky130_fd_sc_hd__and2b_1 _13401_ (.A_N(_06084_),
    .B(_06083_),
    .X(_06090_));
 sky130_fd_sc_hd__xnor2_1 _13402_ (.A(_06068_),
    .B(_06088_),
    .Y(_06091_));
 sky130_fd_sc_hd__nand2_1 _13403_ (.A(_06090_),
    .B(_06091_),
    .Y(_06092_));
 sky130_fd_sc_hd__xnor2_1 _13404_ (.A(_06037_),
    .B(_06057_),
    .Y(_06093_));
 sky130_fd_sc_hd__a21oi_1 _13405_ (.A1(_06089_),
    .A2(_06092_),
    .B1(_06093_),
    .Y(_06094_));
 sky130_fd_sc_hd__inv_2 _13406_ (.A(_06094_),
    .Y(_06095_));
 sky130_fd_sc_hd__or2_1 _13407_ (.A(_06090_),
    .B(_06091_),
    .X(_06096_));
 sky130_fd_sc_hd__or2_1 _13408_ (.A(_06085_),
    .B(_06086_),
    .X(_06097_));
 sky130_fd_sc_hd__and2_1 _13409_ (.A(_06087_),
    .B(_06097_),
    .X(_06098_));
 sky130_fd_sc_hd__nand3_1 _13410_ (.A(_06073_),
    .B(_06074_),
    .C(_06080_),
    .Y(_06099_));
 sky130_fd_sc_hd__a21o_1 _13411_ (.A1(_06073_),
    .A2(_06074_),
    .B1(_06080_),
    .X(_06100_));
 sky130_fd_sc_hd__clkbuf_4 _13412_ (.A(_05631_),
    .X(_06101_));
 sky130_fd_sc_hd__or4_1 _13413_ (.A(_05671_),
    .B(_05629_),
    .C(_05622_),
    .D(_06101_),
    .X(_06102_));
 sky130_fd_sc_hd__a22o_1 _13414_ (.A1(_05699_),
    .A2(_05641_),
    .B1(_05651_),
    .B2(_05612_),
    .X(_06103_));
 sky130_fd_sc_hd__nand4_1 _13415_ (.A(_06028_),
    .B(_05738_),
    .C(_06102_),
    .D(_06103_),
    .Y(_06104_));
 sky130_fd_sc_hd__a22o_1 _13416_ (.A1(_06028_),
    .A2(_05738_),
    .B1(_06102_),
    .B2(_06103_),
    .X(_06105_));
 sky130_fd_sc_hd__xnor2_1 _13417_ (.A(_06077_),
    .B(_06078_),
    .Y(_06106_));
 sky130_fd_sc_hd__nor2_1 _13418_ (.A(_05793_),
    .B(_05635_),
    .Y(_06107_));
 sky130_fd_sc_hd__or3b_1 _13419_ (.A(_05625_),
    .B(_05959_),
    .C_N(_06107_),
    .X(_06108_));
 sky130_fd_sc_hd__a21o_1 _13420_ (.A1(_05525_),
    .A2(_05668_),
    .B1(_06107_),
    .X(_06109_));
 sky130_fd_sc_hd__a21bo_1 _13421_ (.A1(_06007_),
    .A2(_06108_),
    .B1_N(_06109_),
    .X(_06110_));
 sky130_fd_sc_hd__nand2_1 _13422_ (.A(_06106_),
    .B(_06110_),
    .Y(_06111_));
 sky130_fd_sc_hd__nor2_1 _13423_ (.A(_06106_),
    .B(_06110_),
    .Y(_06112_));
 sky130_fd_sc_hd__a31o_1 _13424_ (.A1(_06104_),
    .A2(_06105_),
    .A3(_06111_),
    .B1(_06112_),
    .X(_06113_));
 sky130_fd_sc_hd__and3_1 _13425_ (.A(_06099_),
    .B(_06100_),
    .C(_06113_),
    .X(_06114_));
 sky130_fd_sc_hd__nand2_2 _13426_ (.A(_05618_),
    .B(_05745_),
    .Y(_06115_));
 sky130_fd_sc_hd__nand2_1 _13427_ (.A(_06028_),
    .B(_06115_),
    .Y(_06116_));
 sky130_fd_sc_hd__and2_1 _13428_ (.A(_06102_),
    .B(_06104_),
    .X(_06117_));
 sky130_fd_sc_hd__xnor2_1 _13429_ (.A(_06116_),
    .B(_06117_),
    .Y(_06118_));
 sky130_fd_sc_hd__a21oi_1 _13430_ (.A1(_06099_),
    .A2(_06100_),
    .B1(_06113_),
    .Y(_06119_));
 sky130_fd_sc_hd__nor3_1 _13431_ (.A(_06114_),
    .B(_06118_),
    .C(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__or3_1 _13432_ (.A(_06098_),
    .B(_06114_),
    .C(_06120_),
    .X(_06121_));
 sky130_fd_sc_hd__xnor2_1 _13433_ (.A(_05612_),
    .B(_05525_),
    .Y(_06122_));
 sky130_fd_sc_hd__or4_1 _13434_ (.A(_05793_),
    .B(_05671_),
    .C(_05740_),
    .D(_06122_),
    .X(_06123_));
 sky130_fd_sc_hd__and2_1 _13435_ (.A(_06104_),
    .B(_06105_),
    .X(_06124_));
 sky130_fd_sc_hd__or2b_1 _13436_ (.A(_06112_),
    .B_N(_06111_),
    .X(_06125_));
 sky130_fd_sc_hd__xnor2_1 _13437_ (.A(_06124_),
    .B(_06125_),
    .Y(_06126_));
 sky130_fd_sc_hd__inv_2 _13438_ (.A(_06007_),
    .Y(_06127_));
 sky130_fd_sc_hd__nand2_1 _13439_ (.A(_06108_),
    .B(_06109_),
    .Y(_06128_));
 sky130_fd_sc_hd__nand2_1 _13440_ (.A(_05488_),
    .B(_05625_),
    .Y(_06129_));
 sky130_fd_sc_hd__o211a_1 _13441_ (.A1(_05629_),
    .A2(_06129_),
    .B1(_06109_),
    .C1(_06108_),
    .X(_06130_));
 sky130_fd_sc_hd__a41o_1 _13442_ (.A1(_06028_),
    .A2(_05612_),
    .A3(_05625_),
    .A4(_05715_),
    .B1(_06130_),
    .X(_06131_));
 sky130_fd_sc_hd__a2bb2o_1 _13443_ (.A1_N(_06122_),
    .A2_N(_05671_),
    .B1(_06028_),
    .B2(_05641_),
    .X(_06132_));
 sky130_fd_sc_hd__and2_1 _13444_ (.A(_06123_),
    .B(_06132_),
    .X(_06133_));
 sky130_fd_sc_hd__a32o_1 _13445_ (.A1(_06127_),
    .A2(_06128_),
    .A3(_06129_),
    .B1(_06131_),
    .B2(_06133_),
    .X(_06134_));
 sky130_fd_sc_hd__nand2_1 _13446_ (.A(_06126_),
    .B(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__nor2_1 _13447_ (.A(_06126_),
    .B(_06134_),
    .Y(_06136_));
 sky130_fd_sc_hd__clkbuf_4 _13448_ (.A(_05793_),
    .X(_06137_));
 sky130_fd_sc_hd__a211o_1 _13449_ (.A1(_06133_),
    .A2(_06131_),
    .B1(_06137_),
    .C1(_06122_),
    .X(_06138_));
 sky130_fd_sc_hd__nor2_1 _13450_ (.A(_06133_),
    .B(_06131_),
    .Y(_06139_));
 sky130_fd_sc_hd__or3_1 _13451_ (.A(_06136_),
    .B(_06138_),
    .C(_06139_),
    .X(_06140_));
 sky130_fd_sc_hd__o21a_1 _13452_ (.A1(_06114_),
    .A2(_06119_),
    .B1(_06118_),
    .X(_06141_));
 sky130_fd_sc_hd__a31o_1 _13453_ (.A1(_06123_),
    .A2(_06135_),
    .A3(_06140_),
    .B1(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__o21ai_1 _13454_ (.A1(_06114_),
    .A2(_06120_),
    .B1(_06098_),
    .Y(_06143_));
 sky130_fd_sc_hd__o221ai_1 _13455_ (.A1(_06116_),
    .A2(_06117_),
    .B1(_06120_),
    .B2(_06142_),
    .C1(_06143_),
    .Y(_06144_));
 sky130_fd_sc_hd__and4_1 _13456_ (.A(_06092_),
    .B(_06096_),
    .C(_06121_),
    .D(_06144_),
    .X(_06145_));
 sky130_fd_sc_hd__nand3_1 _13457_ (.A(_06093_),
    .B(_06089_),
    .C(_06092_),
    .Y(_06146_));
 sky130_fd_sc_hd__and3_1 _13458_ (.A(_06095_),
    .B(_06145_),
    .C(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__and4bb_1 _13459_ (.A_N(_06066_),
    .B_N(_06067_),
    .C(_06147_),
    .D(_06095_),
    .X(_06148_));
 sky130_fd_sc_hd__a211o_1 _13460_ (.A1(_06064_),
    .A2(_06060_),
    .B1(_06095_),
    .C1(_06066_),
    .X(_06149_));
 sky130_fd_sc_hd__or3b_1 _13461_ (.A(_06026_),
    .B(_06065_),
    .C_N(_06149_),
    .X(_06150_));
 sky130_fd_sc_hd__a21o_1 _13462_ (.A1(_06060_),
    .A2(_06063_),
    .B1(_06064_),
    .X(_06151_));
 sky130_fd_sc_hd__xnor2_1 _13463_ (.A(_05981_),
    .B(_06022_),
    .Y(_06152_));
 sky130_fd_sc_hd__a21o_1 _13464_ (.A1(_06151_),
    .A2(_06149_),
    .B1(_06152_),
    .X(_06153_));
 sky130_fd_sc_hd__nor2_1 _13465_ (.A(_06152_),
    .B(_06149_),
    .Y(_06154_));
 sky130_fd_sc_hd__a31o_1 _13466_ (.A1(_06148_),
    .A2(_06150_),
    .A3(_06153_),
    .B1(_06154_),
    .X(_06155_));
 sky130_fd_sc_hd__a21oi_1 _13467_ (.A1(_06026_),
    .A2(_06065_),
    .B1(_06023_),
    .Y(_06156_));
 sky130_fd_sc_hd__xnor2_1 _13468_ (.A(_06024_),
    .B(_06156_),
    .Y(_06157_));
 sky130_fd_sc_hd__a32o_1 _13469_ (.A1(_06024_),
    .A2(_06026_),
    .A3(_06065_),
    .B1(_06155_),
    .B2(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__nor3_1 _13470_ (.A(_05978_),
    .B(_05979_),
    .C(_06025_),
    .Y(_06159_));
 sky130_fd_sc_hd__a211oi_1 _13471_ (.A1(_05979_),
    .A2(_06025_),
    .B1(_06159_),
    .C1(_05980_),
    .Y(_06160_));
 sky130_fd_sc_hd__a22o_1 _13472_ (.A1(_05979_),
    .A2(_06025_),
    .B1(_06158_),
    .B2(_06160_),
    .X(_06161_));
 sky130_fd_sc_hd__nor2_1 _13473_ (.A(_05934_),
    .B(_05980_),
    .Y(_06162_));
 sky130_fd_sc_hd__xnor2_1 _13474_ (.A(_05881_),
    .B(_06162_),
    .Y(_06163_));
 sky130_fd_sc_hd__a22o_1 _13475_ (.A1(_05881_),
    .A2(_05980_),
    .B1(_06161_),
    .B2(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__xor2_1 _13476_ (.A(_05936_),
    .B(_06164_),
    .X(_06165_));
 sky130_fd_sc_hd__xor2_1 _13477_ (.A(_06161_),
    .B(_06163_),
    .X(_06166_));
 sky130_fd_sc_hd__xor2_1 _13478_ (.A(_06158_),
    .B(_06160_),
    .X(_06167_));
 sky130_fd_sc_hd__xnor2_1 _13479_ (.A(_06155_),
    .B(_06157_),
    .Y(_06168_));
 sky130_fd_sc_hd__and3_1 _13480_ (.A(_06148_),
    .B(_06150_),
    .C(_06153_),
    .X(_06169_));
 sky130_fd_sc_hd__a21oi_1 _13481_ (.A1(_06150_),
    .A2(_06153_),
    .B1(_06148_),
    .Y(_06170_));
 sky130_fd_sc_hd__or2_1 _13482_ (.A(_06169_),
    .B(_06170_),
    .X(_06171_));
 sky130_fd_sc_hd__buf_2 _13483_ (.A(_06171_),
    .X(_06172_));
 sky130_fd_sc_hd__nand2_1 _13484_ (.A(_06168_),
    .B(_06172_),
    .Y(_06173_));
 sky130_fd_sc_hd__and2_1 _13485_ (.A(_06167_),
    .B(_06173_),
    .X(_06174_));
 sky130_fd_sc_hd__or2_1 _13486_ (.A(_06166_),
    .B(_06174_),
    .X(_06175_));
 sky130_fd_sc_hd__or2_2 _13487_ (.A(_06165_),
    .B(_06175_),
    .X(_06176_));
 sky130_fd_sc_hd__nand2_1 _13488_ (.A(_05839_),
    .B(_05878_),
    .Y(_06177_));
 sky130_fd_sc_hd__and2b_1 _13489_ (.A_N(_05877_),
    .B(_05842_),
    .X(_06178_));
 sky130_fd_sc_hd__or2b_1 _13490_ (.A(_05876_),
    .B_N(_05874_),
    .X(_06179_));
 sky130_fd_sc_hd__and2b_1 _13491_ (.A_N(_05856_),
    .B(_05870_),
    .X(_06180_));
 sky130_fd_sc_hd__a21o_1 _13492_ (.A1(_05756_),
    .A2(_05855_),
    .B1(_06180_),
    .X(_06181_));
 sky130_fd_sc_hd__and3_1 _13493_ (.A(_05401_),
    .B(_05738_),
    .C(_05854_),
    .X(_06182_));
 sky130_fd_sc_hd__inv_2 _13494_ (.A(_05847_),
    .Y(_06183_));
 sky130_fd_sc_hd__o21ba_1 _13495_ (.A1(_06183_),
    .A2(_05850_),
    .B1_N(_05849_),
    .X(_06184_));
 sky130_fd_sc_hd__a21oi_1 _13496_ (.A1(_05401_),
    .A2(_06115_),
    .B1(_05848_),
    .Y(_06185_));
 sky130_fd_sc_hd__and2_1 _13497_ (.A(_06115_),
    .B(_05848_),
    .X(_06186_));
 sky130_fd_sc_hd__nor4_2 _13498_ (.A(_05621_),
    .B(_05610_),
    .C(_06185_),
    .D(_06186_),
    .Y(_06187_));
 sky130_fd_sc_hd__o22a_1 _13499_ (.A1(_05621_),
    .A2(_05610_),
    .B1(_06185_),
    .B2(_06186_),
    .X(_06188_));
 sky130_fd_sc_hd__nor2_1 _13500_ (.A(_06187_),
    .B(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__xnor2_1 _13501_ (.A(_06184_),
    .B(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__nand2_1 _13502_ (.A(_06182_),
    .B(_06190_),
    .Y(_06191_));
 sky130_fd_sc_hd__or2_1 _13503_ (.A(_06182_),
    .B(_06190_),
    .X(_06192_));
 sky130_fd_sc_hd__and2_1 _13504_ (.A(_06191_),
    .B(_06192_),
    .X(_06193_));
 sky130_fd_sc_hd__or2b_1 _13505_ (.A(_05853_),
    .B_N(_05846_),
    .X(_06194_));
 sky130_fd_sc_hd__a21bo_1 _13506_ (.A1(_05739_),
    .A2(_05852_),
    .B1_N(_06194_),
    .X(_06195_));
 sky130_fd_sc_hd__and3_1 _13507_ (.A(_05692_),
    .B(_05722_),
    .C(_05772_),
    .X(_06196_));
 sky130_fd_sc_hd__and2b_1 _13508_ (.A_N(_05862_),
    .B(_05864_),
    .X(_06197_));
 sky130_fd_sc_hd__nand2_1 _13509_ (.A(_05692_),
    .B(_05722_),
    .Y(_06198_));
 sky130_fd_sc_hd__nor2_1 _13510_ (.A(_05608_),
    .B(_05767_),
    .Y(_06199_));
 sky130_fd_sc_hd__xnor2_1 _13511_ (.A(_06198_),
    .B(_06199_),
    .Y(_06200_));
 sky130_fd_sc_hd__and3_1 _13512_ (.A(_05553_),
    .B(_05701_),
    .C(_06200_),
    .X(_06201_));
 sky130_fd_sc_hd__a21oi_1 _13513_ (.A1(_05553_),
    .A2(_05701_),
    .B1(_06200_),
    .Y(_06202_));
 sky130_fd_sc_hd__nor2_1 _13514_ (.A(_06201_),
    .B(_06202_),
    .Y(_06203_));
 sky130_fd_sc_hd__o21ai_1 _13515_ (.A1(_06196_),
    .A2(_06197_),
    .B1(_06203_),
    .Y(_06204_));
 sky130_fd_sc_hd__or3_1 _13516_ (.A(_06196_),
    .B(_06197_),
    .C(_06203_),
    .X(_06205_));
 sky130_fd_sc_hd__and2_1 _13517_ (.A(_06204_),
    .B(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__xnor2_1 _13518_ (.A(_06195_),
    .B(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__xor2_1 _13519_ (.A(_05866_),
    .B(_06207_),
    .X(_06208_));
 sky130_fd_sc_hd__xnor2_1 _13520_ (.A(_06193_),
    .B(_06208_),
    .Y(_06209_));
 sky130_fd_sc_hd__xnor2_1 _13521_ (.A(_06181_),
    .B(_06209_),
    .Y(_06210_));
 sky130_fd_sc_hd__nor2_1 _13522_ (.A(_05775_),
    .B(_05869_),
    .Y(_06211_));
 sky130_fd_sc_hd__a21oi_1 _13523_ (.A1(_05858_),
    .A2(_05868_),
    .B1(_06211_),
    .Y(_06212_));
 sky130_fd_sc_hd__xor2_1 _13524_ (.A(_06210_),
    .B(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__a21oi_2 _13525_ (.A1(_05872_),
    .A2(_06179_),
    .B1(_06213_),
    .Y(_06214_));
 sky130_fd_sc_hd__and3_1 _13526_ (.A(_05872_),
    .B(_06179_),
    .C(_06213_),
    .X(_06215_));
 sky130_fd_sc_hd__nor2_1 _13527_ (.A(_06214_),
    .B(_06215_),
    .Y(_06216_));
 sky130_fd_sc_hd__xor2_1 _13528_ (.A(_06178_),
    .B(_06216_),
    .X(_06217_));
 sky130_fd_sc_hd__xnor2_1 _13529_ (.A(_06177_),
    .B(_06217_),
    .Y(_06218_));
 sky130_fd_sc_hd__and2_1 _13530_ (.A(_05879_),
    .B(_05935_),
    .X(_06219_));
 sky130_fd_sc_hd__a21o_1 _13531_ (.A1(_05936_),
    .A2(_06164_),
    .B1(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__xor2_1 _13532_ (.A(_06218_),
    .B(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__or2_2 _13533_ (.A(_06176_),
    .B(_06221_),
    .X(_06222_));
 sky130_fd_sc_hd__and3_1 _13534_ (.A(_05839_),
    .B(_05878_),
    .C(_06217_),
    .X(_06223_));
 sky130_fd_sc_hd__a21o_1 _13535_ (.A1(_06218_),
    .A2(_06220_),
    .B1(_06223_),
    .X(_06224_));
 sky130_fd_sc_hd__and2_1 _13536_ (.A(_06178_),
    .B(_06216_),
    .X(_06225_));
 sky130_fd_sc_hd__or2b_1 _13537_ (.A(_06209_),
    .B_N(_06181_),
    .X(_06226_));
 sky130_fd_sc_hd__or2b_1 _13538_ (.A(_06212_),
    .B_N(_06210_),
    .X(_06227_));
 sky130_fd_sc_hd__nand2_1 _13539_ (.A(_06226_),
    .B(_06227_),
    .Y(_06228_));
 sky130_fd_sc_hd__a21bo_1 _13540_ (.A1(_06193_),
    .A2(_06208_),
    .B1_N(_06191_),
    .X(_06229_));
 sky130_fd_sc_hd__inv_2 _13541_ (.A(_05610_),
    .Y(_06230_));
 sky130_fd_sc_hd__nand2_1 _13542_ (.A(_06230_),
    .B(_05848_),
    .Y(_06231_));
 sky130_fd_sc_hd__o21ai_1 _13543_ (.A1(_05624_),
    .A2(_05610_),
    .B1(_05749_),
    .Y(_06232_));
 sky130_fd_sc_hd__and2_1 _13544_ (.A(_06231_),
    .B(_06232_),
    .X(_06233_));
 sky130_fd_sc_hd__o21a_1 _13545_ (.A1(_06186_),
    .A2(_06187_),
    .B1(_06233_),
    .X(_06234_));
 sky130_fd_sc_hd__nor3_1 _13546_ (.A(_06186_),
    .B(_06187_),
    .C(_06233_),
    .Y(_06235_));
 sky130_fd_sc_hd__nor2_1 _13547_ (.A(_06234_),
    .B(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__or3_1 _13548_ (.A(_06184_),
    .B(_06187_),
    .C(_06188_),
    .X(_06237_));
 sky130_fd_sc_hd__and3_1 _13549_ (.A(_05692_),
    .B(_05722_),
    .C(_06199_),
    .X(_06238_));
 sky130_fd_sc_hd__or4_1 _13550_ (.A(_05433_),
    .B(_05608_),
    .C(_05611_),
    .D(_05583_),
    .X(_06239_));
 sky130_fd_sc_hd__a22o_1 _13551_ (.A1(_05645_),
    .A2(_05624_),
    .B1(_05701_),
    .B2(_05692_),
    .X(_06240_));
 sky130_fd_sc_hd__and2_1 _13552_ (.A(_06239_),
    .B(_06240_),
    .X(_06241_));
 sky130_fd_sc_hd__o21ai_2 _13553_ (.A1(_06238_),
    .A2(_06201_),
    .B1(_06241_),
    .Y(_06242_));
 sky130_fd_sc_hd__or3_1 _13554_ (.A(_06238_),
    .B(_06201_),
    .C(_06241_),
    .X(_06243_));
 sky130_fd_sc_hd__and2_1 _13555_ (.A(_06242_),
    .B(_06243_),
    .X(_06244_));
 sky130_fd_sc_hd__xor2_1 _13556_ (.A(_06237_),
    .B(_06244_),
    .X(_06245_));
 sky130_fd_sc_hd__xor2_1 _13557_ (.A(_06204_),
    .B(_06245_),
    .X(_06246_));
 sky130_fd_sc_hd__nand2_1 _13558_ (.A(_06236_),
    .B(_06246_),
    .Y(_06247_));
 sky130_fd_sc_hd__or2_1 _13559_ (.A(_06236_),
    .B(_06246_),
    .X(_06248_));
 sky130_fd_sc_hd__nand2_1 _13560_ (.A(_06247_),
    .B(_06248_),
    .Y(_06249_));
 sky130_fd_sc_hd__xnor2_1 _13561_ (.A(_06229_),
    .B(_06249_),
    .Y(_06250_));
 sky130_fd_sc_hd__nor2_1 _13562_ (.A(_05866_),
    .B(_06207_),
    .Y(_06251_));
 sky130_fd_sc_hd__a21oi_1 _13563_ (.A1(_06195_),
    .A2(_06206_),
    .B1(_06251_),
    .Y(_06252_));
 sky130_fd_sc_hd__xor2_1 _13564_ (.A(_06250_),
    .B(_06252_),
    .X(_06253_));
 sky130_fd_sc_hd__xnor2_2 _13565_ (.A(_06228_),
    .B(_06253_),
    .Y(_06254_));
 sky130_fd_sc_hd__xor2_1 _13566_ (.A(_06214_),
    .B(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__and2_1 _13567_ (.A(_06225_),
    .B(_06255_),
    .X(_06256_));
 sky130_fd_sc_hd__nor2_1 _13568_ (.A(_06225_),
    .B(_06255_),
    .Y(_06257_));
 sky130_fd_sc_hd__nor2_1 _13569_ (.A(_06256_),
    .B(_06257_),
    .Y(_06258_));
 sky130_fd_sc_hd__xor2_2 _13570_ (.A(_06224_),
    .B(_06258_),
    .X(_06259_));
 sky130_fd_sc_hd__nor2_2 _13571_ (.A(_06222_),
    .B(_06259_),
    .Y(_06260_));
 sky130_fd_sc_hd__a21o_1 _13572_ (.A1(_06224_),
    .A2(_06258_),
    .B1(_06256_),
    .X(_06261_));
 sky130_fd_sc_hd__nand2_2 _13573_ (.A(_06214_),
    .B(_06254_),
    .Y(_06262_));
 sky130_fd_sc_hd__and2b_1 _13574_ (.A_N(_06253_),
    .B(_06228_),
    .X(_06263_));
 sky130_fd_sc_hd__and2b_1 _13575_ (.A_N(_06252_),
    .B(_06250_),
    .X(_06264_));
 sky130_fd_sc_hd__a31o_1 _13576_ (.A1(_06229_),
    .A2(_06247_),
    .A3(_06248_),
    .B1(_06264_),
    .X(_06265_));
 sky130_fd_sc_hd__clkbuf_4 _13577_ (.A(_05610_),
    .X(_06266_));
 sky130_fd_sc_hd__or3_1 _13578_ (.A(_05434_),
    .B(_06266_),
    .C(_05848_),
    .X(_06267_));
 sky130_fd_sc_hd__nand2_1 _13579_ (.A(_05645_),
    .B(_05701_),
    .Y(_06268_));
 sky130_fd_sc_hd__nand2_1 _13580_ (.A(_05621_),
    .B(_05624_),
    .Y(_06269_));
 sky130_fd_sc_hd__and3_1 _13581_ (.A(_06183_),
    .B(_05702_),
    .C(_06269_),
    .X(_06270_));
 sky130_fd_sc_hd__xnor2_1 _13582_ (.A(_06268_),
    .B(_06270_),
    .Y(_06271_));
 sky130_fd_sc_hd__o21a_1 _13583_ (.A1(_05606_),
    .A2(_06271_),
    .B1(_06239_),
    .X(_06272_));
 sky130_fd_sc_hd__nand2_1 _13584_ (.A(_06234_),
    .B(_06272_),
    .Y(_06273_));
 sky130_fd_sc_hd__or2_1 _13585_ (.A(_06234_),
    .B(_06272_),
    .X(_06274_));
 sky130_fd_sc_hd__nand2_1 _13586_ (.A(_06273_),
    .B(_06274_),
    .Y(_06275_));
 sky130_fd_sc_hd__xnor2_1 _13587_ (.A(_06242_),
    .B(_06275_),
    .Y(_06276_));
 sky130_fd_sc_hd__nor2_1 _13588_ (.A(_06267_),
    .B(_06276_),
    .Y(_06277_));
 sky130_fd_sc_hd__and2_1 _13589_ (.A(_06267_),
    .B(_06276_),
    .X(_06278_));
 sky130_fd_sc_hd__nor2_1 _13590_ (.A(_06277_),
    .B(_06278_),
    .Y(_06279_));
 sky130_fd_sc_hd__xnor2_1 _13591_ (.A(_06247_),
    .B(_06279_),
    .Y(_06280_));
 sky130_fd_sc_hd__and2b_1 _13592_ (.A_N(_06237_),
    .B(_06244_),
    .X(_06281_));
 sky130_fd_sc_hd__o21bai_1 _13593_ (.A1(_06204_),
    .A2(_06245_),
    .B1_N(_06281_),
    .Y(_06282_));
 sky130_fd_sc_hd__xnor2_1 _13594_ (.A(_06280_),
    .B(_06282_),
    .Y(_06283_));
 sky130_fd_sc_hd__xnor2_1 _13595_ (.A(_06265_),
    .B(_06283_),
    .Y(_06284_));
 sky130_fd_sc_hd__and2_1 _13596_ (.A(_06263_),
    .B(_06284_),
    .X(_06285_));
 sky130_fd_sc_hd__nor2_1 _13597_ (.A(_06263_),
    .B(_06284_),
    .Y(_06286_));
 sky130_fd_sc_hd__nor2_2 _13598_ (.A(_06285_),
    .B(_06286_),
    .Y(_06287_));
 sky130_fd_sc_hd__xnor2_4 _13599_ (.A(_06262_),
    .B(_06287_),
    .Y(_06288_));
 sky130_fd_sc_hd__xnor2_4 _13600_ (.A(_06261_),
    .B(_06288_),
    .Y(_06289_));
 sky130_fd_sc_hd__and2_1 _13601_ (.A(_06224_),
    .B(_06258_),
    .X(_06290_));
 sky130_fd_sc_hd__and2b_1 _13602_ (.A_N(_06283_),
    .B(_06265_),
    .X(_06291_));
 sky130_fd_sc_hd__a32o_1 _13603_ (.A1(_06236_),
    .A2(_06246_),
    .A3(_06279_),
    .B1(_06280_),
    .B2(_06282_),
    .X(_06292_));
 sky130_fd_sc_hd__or2_1 _13604_ (.A(_05434_),
    .B(_05847_),
    .X(_06293_));
 sky130_fd_sc_hd__a32o_1 _13605_ (.A1(_05645_),
    .A2(_05701_),
    .A3(_06270_),
    .B1(_06293_),
    .B2(_05703_),
    .X(_06294_));
 sky130_fd_sc_hd__xnor2_1 _13606_ (.A(_06231_),
    .B(_06294_),
    .Y(_06295_));
 sky130_fd_sc_hd__nand2_1 _13607_ (.A(_06239_),
    .B(_06295_),
    .Y(_06296_));
 sky130_fd_sc_hd__o221a_1 _13608_ (.A1(_06242_),
    .A2(_06275_),
    .B1(_06277_),
    .B2(_06296_),
    .C1(_06273_),
    .X(_06297_));
 sky130_fd_sc_hd__a21bo_1 _13609_ (.A1(_06277_),
    .A2(_06296_),
    .B1_N(_06297_),
    .X(_06298_));
 sky130_fd_sc_hd__xnor2_1 _13610_ (.A(_06292_),
    .B(_06298_),
    .Y(_06299_));
 sky130_fd_sc_hd__xnor2_1 _13611_ (.A(_06291_),
    .B(_06299_),
    .Y(_06300_));
 sky130_fd_sc_hd__a21o_1 _13612_ (.A1(_06214_),
    .A2(_06254_),
    .B1(_06256_),
    .X(_06301_));
 sky130_fd_sc_hd__a21o_1 _13613_ (.A1(_06287_),
    .A2(_06301_),
    .B1(_06285_),
    .X(_06302_));
 sky130_fd_sc_hd__a211oi_2 _13614_ (.A1(_06290_),
    .A2(_06288_),
    .B1(_06300_),
    .C1(_06302_),
    .Y(_06303_));
 sky130_fd_sc_hd__a21oi_1 _13615_ (.A1(_06260_),
    .A2(_06289_),
    .B1(_06303_),
    .Y(_06304_));
 sky130_fd_sc_hd__buf_2 _13616_ (.A(_06304_),
    .X(_06305_));
 sky130_fd_sc_hd__buf_2 _13617_ (.A(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__nor2_1 _13618_ (.A(_05606_),
    .B(_06306_),
    .Y(_06307_));
 sky130_fd_sc_hd__o21a_1 _13619_ (.A1(_05722_),
    .A2(_05818_),
    .B1(_06306_),
    .X(_06308_));
 sky130_fd_sc_hd__nand2_1 _13620_ (.A(_06230_),
    .B(_06306_),
    .Y(_06309_));
 sky130_fd_sc_hd__buf_2 _13621_ (.A(_05746_),
    .X(_06310_));
 sky130_fd_sc_hd__nor2_1 _13622_ (.A(_05434_),
    .B(_06306_),
    .Y(_06311_));
 sky130_fd_sc_hd__inv_2 _13623_ (.A(_06311_),
    .Y(_06312_));
 sky130_fd_sc_hd__clkbuf_4 _13624_ (.A(_05749_),
    .X(_06313_));
 sky130_fd_sc_hd__or2b_1 _13625_ (.A(_06313_),
    .B_N(_06305_),
    .X(_06314_));
 sky130_fd_sc_hd__o21a_1 _13626_ (.A1(_06310_),
    .A2(_06312_),
    .B1(_06314_),
    .X(_06315_));
 sky130_fd_sc_hd__nor2_1 _13627_ (.A(_06309_),
    .B(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__buf_2 _13628_ (.A(_05728_),
    .X(_06317_));
 sky130_fd_sc_hd__nand2_1 _13629_ (.A(_05818_),
    .B(_06306_),
    .Y(_06318_));
 sky130_fd_sc_hd__or2_1 _13630_ (.A(_06317_),
    .B(_06318_),
    .X(_06319_));
 sky130_fd_sc_hd__xor2_4 _13631_ (.A(_06260_),
    .B(_06289_),
    .X(_06320_));
 sky130_fd_sc_hd__buf_2 _13632_ (.A(_06320_),
    .X(_06321_));
 sky130_fd_sc_hd__and3_1 _13633_ (.A(_05701_),
    .B(_06319_),
    .C(_06321_),
    .X(_06322_));
 sky130_fd_sc_hd__and2_1 _13634_ (.A(_06316_),
    .B(_06322_),
    .X(_06323_));
 sky130_fd_sc_hd__or2_1 _13635_ (.A(_06310_),
    .B(_06314_),
    .X(_06324_));
 sky130_fd_sc_hd__and2_1 _13636_ (.A(_06115_),
    .B(_06305_),
    .X(_06325_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13637_ (.A(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__xor2_2 _13638_ (.A(_06314_),
    .B(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__or2_1 _13639_ (.A(_06309_),
    .B(_06327_),
    .X(_06328_));
 sky130_fd_sc_hd__a21o_1 _13640_ (.A1(_06324_),
    .A2(_06328_),
    .B1(_06316_),
    .X(_06329_));
 sky130_fd_sc_hd__xnor2_2 _13641_ (.A(_06222_),
    .B(_06259_),
    .Y(_06330_));
 sky130_fd_sc_hd__buf_2 _13642_ (.A(_06330_),
    .X(_06331_));
 sky130_fd_sc_hd__nor2_1 _13643_ (.A(_05861_),
    .B(_06331_),
    .Y(_06332_));
 sky130_fd_sc_hd__and2_1 _13644_ (.A(_05722_),
    .B(_06321_),
    .X(_06333_));
 sky130_fd_sc_hd__mux2_1 _13645_ (.A0(_06317_),
    .A1(_06333_),
    .S(_06318_),
    .X(_06334_));
 sky130_fd_sc_hd__a21boi_1 _13646_ (.A1(_06332_),
    .A2(_06334_),
    .B1_N(_06319_),
    .Y(_06335_));
 sky130_fd_sc_hd__nand2_1 _13647_ (.A(_06308_),
    .B(_06322_),
    .Y(_06336_));
 sky130_fd_sc_hd__and3_1 _13648_ (.A(_06306_),
    .B(_06335_),
    .C(_06336_),
    .X(_06337_));
 sky130_fd_sc_hd__inv_2 _13649_ (.A(_06337_),
    .Y(_06338_));
 sky130_fd_sc_hd__xnor2_1 _13650_ (.A(_06332_),
    .B(_06334_),
    .Y(_06339_));
 sky130_fd_sc_hd__nor2_1 _13651_ (.A(_05767_),
    .B(_06331_),
    .Y(_06340_));
 sky130_fd_sc_hd__nand2_1 _13652_ (.A(_06176_),
    .B(_06221_),
    .Y(_06341_));
 sky130_fd_sc_hd__nand2_1 _13653_ (.A(_06222_),
    .B(_06341_),
    .Y(_06342_));
 sky130_fd_sc_hd__clkbuf_4 _13654_ (.A(_06342_),
    .X(_06343_));
 sky130_fd_sc_hd__nor2_1 _13655_ (.A(_05861_),
    .B(_06343_),
    .Y(_06344_));
 sky130_fd_sc_hd__o2bb2a_1 _13656_ (.A1_N(_05818_),
    .A2_N(_06321_),
    .B1(_06331_),
    .B2(_06317_),
    .X(_06345_));
 sky130_fd_sc_hd__a21oi_2 _13657_ (.A1(_06333_),
    .A2(_06340_),
    .B1(_06345_),
    .Y(_06346_));
 sky130_fd_sc_hd__a22oi_1 _13658_ (.A1(_06333_),
    .A2(_06340_),
    .B1(_06344_),
    .B2(_06346_),
    .Y(_06347_));
 sky130_fd_sc_hd__or2_1 _13659_ (.A(_06339_),
    .B(_06347_),
    .X(_06348_));
 sky130_fd_sc_hd__xnor2_1 _13660_ (.A(_06329_),
    .B(_06337_),
    .Y(_06349_));
 sky130_fd_sc_hd__or2b_1 _13661_ (.A(_06348_),
    .B_N(_06349_),
    .X(_06350_));
 sky130_fd_sc_hd__o21ai_1 _13662_ (.A1(_06329_),
    .A2(_06338_),
    .B1(_06350_),
    .Y(_06351_));
 sky130_fd_sc_hd__o21a_1 _13663_ (.A1(_06313_),
    .A2(_06306_),
    .B1(_06309_),
    .X(_06352_));
 sky130_fd_sc_hd__a21o_1 _13664_ (.A1(_05401_),
    .A2(_06352_),
    .B1(_06316_),
    .X(_06353_));
 sky130_fd_sc_hd__xnor2_1 _13665_ (.A(_06348_),
    .B(_06349_),
    .Y(_06354_));
 sky130_fd_sc_hd__and2b_1 _13666_ (.A_N(_06353_),
    .B(_06354_),
    .X(_06355_));
 sky130_fd_sc_hd__nor2_1 _13667_ (.A(_06316_),
    .B(_06322_),
    .Y(_06356_));
 sky130_fd_sc_hd__o21ai_1 _13668_ (.A1(_06323_),
    .A2(_06356_),
    .B1(_06335_),
    .Y(_06357_));
 sky130_fd_sc_hd__or3_1 _13669_ (.A(_06323_),
    .B(_06335_),
    .C(_06356_),
    .X(_06358_));
 sky130_fd_sc_hd__o2bb2a_1 _13670_ (.A1_N(_06357_),
    .A2_N(_06358_),
    .B1(_06266_),
    .B2(_06312_),
    .X(_06359_));
 sky130_fd_sc_hd__nor2_1 _13671_ (.A(_06355_),
    .B(_06359_),
    .Y(_06360_));
 sky130_fd_sc_hd__a21oi_1 _13672_ (.A1(_06351_),
    .A2(_06360_),
    .B1(_06355_),
    .Y(_06361_));
 sky130_fd_sc_hd__o21a_1 _13673_ (.A1(_05722_),
    .A2(_06306_),
    .B1(_06318_),
    .X(_06362_));
 sky130_fd_sc_hd__o21ba_1 _13674_ (.A1(_06316_),
    .A2(_06362_),
    .B1_N(_06323_),
    .X(_06363_));
 sky130_fd_sc_hd__and2b_1 _13675_ (.A_N(_06361_),
    .B(_06363_),
    .X(_06364_));
 sky130_fd_sc_hd__nor2_1 _13676_ (.A(_05722_),
    .B(_06306_),
    .Y(_06365_));
 sky130_fd_sc_hd__o21ai_1 _13677_ (.A1(_06308_),
    .A2(_06365_),
    .B1(_06319_),
    .Y(_06366_));
 sky130_fd_sc_hd__o21a_1 _13678_ (.A1(_06323_),
    .A2(_06364_),
    .B1(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__nor4_4 _13679_ (.A(_05434_),
    .B(_06307_),
    .C(_06308_),
    .D(_06367_),
    .Y(_06368_));
 sky130_fd_sc_hd__or3_1 _13680_ (.A(_06366_),
    .B(_06323_),
    .C(_06364_),
    .X(_06369_));
 sky130_fd_sc_hd__and2b_1 _13681_ (.A_N(_06367_),
    .B(_06369_),
    .X(_06370_));
 sky130_fd_sc_hd__inv_2 _13682_ (.A(_06370_),
    .Y(_06371_));
 sky130_fd_sc_hd__xnor2_1 _13683_ (.A(_06351_),
    .B(_06360_),
    .Y(_06372_));
 sky130_fd_sc_hd__nand2_1 _13684_ (.A(_06309_),
    .B(_06315_),
    .Y(_06373_));
 sky130_fd_sc_hd__a21oi_1 _13685_ (.A1(_06329_),
    .A2(_06373_),
    .B1(_05434_),
    .Y(_06374_));
 sky130_fd_sc_hd__nand2_1 _13686_ (.A(_06309_),
    .B(_06327_),
    .Y(_06375_));
 sky130_fd_sc_hd__nand2_1 _13687_ (.A(_06328_),
    .B(_06375_),
    .Y(_06376_));
 sky130_fd_sc_hd__inv_2 _13688_ (.A(_06327_),
    .Y(_06377_));
 sky130_fd_sc_hd__and2_1 _13689_ (.A(_06230_),
    .B(_06321_),
    .X(_06378_));
 sky130_fd_sc_hd__a21boi_1 _13690_ (.A1(_06377_),
    .A2(_06378_),
    .B1_N(_06324_),
    .Y(_06379_));
 sky130_fd_sc_hd__nor2_1 _13691_ (.A(_06376_),
    .B(_06379_),
    .Y(_06380_));
 sky130_fd_sc_hd__nand2_1 _13692_ (.A(_06339_),
    .B(_06347_),
    .Y(_06381_));
 sky130_fd_sc_hd__and2_1 _13693_ (.A(_06348_),
    .B(_06381_),
    .X(_06382_));
 sky130_fd_sc_hd__and2_1 _13694_ (.A(_06380_),
    .B(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__nor2_1 _13695_ (.A(_06380_),
    .B(_06382_),
    .Y(_06384_));
 sky130_fd_sc_hd__xnor2_2 _13696_ (.A(_06344_),
    .B(_06346_),
    .Y(_06385_));
 sky130_fd_sc_hd__or2_1 _13697_ (.A(_05767_),
    .B(_06331_),
    .X(_06386_));
 sky130_fd_sc_hd__nand2_1 _13698_ (.A(_06165_),
    .B(_06175_),
    .Y(_06387_));
 sky130_fd_sc_hd__nand2_2 _13699_ (.A(_06176_),
    .B(_06387_),
    .Y(_06388_));
 sky130_fd_sc_hd__clkbuf_4 _13700_ (.A(_06388_),
    .X(_06389_));
 sky130_fd_sc_hd__nor2_1 _13701_ (.A(_06317_),
    .B(_06343_),
    .Y(_06390_));
 sky130_fd_sc_hd__xnor2_1 _13702_ (.A(_06386_),
    .B(_06390_),
    .Y(_06391_));
 sky130_fd_sc_hd__or3b_1 _13703_ (.A(_05861_),
    .B(_06389_),
    .C_N(_06391_),
    .X(_06392_));
 sky130_fd_sc_hd__o31a_1 _13704_ (.A1(_06317_),
    .A2(_06386_),
    .A3(_06343_),
    .B1(_06392_),
    .X(_06393_));
 sky130_fd_sc_hd__o22a_1 _13705_ (.A1(_06383_),
    .A2(_06384_),
    .B1(_06385_),
    .B2(_06393_),
    .X(_06394_));
 sky130_fd_sc_hd__nor2_1 _13706_ (.A(_06374_),
    .B(_06394_),
    .Y(_06395_));
 sky130_fd_sc_hd__xnor2_1 _13707_ (.A(_06353_),
    .B(_06354_),
    .Y(_06396_));
 sky130_fd_sc_hd__xor2_1 _13708_ (.A(_06395_),
    .B(_06396_),
    .X(_06397_));
 sky130_fd_sc_hd__and2_1 _13709_ (.A(_06383_),
    .B(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__a21oi_1 _13710_ (.A1(_06395_),
    .A2(_06396_),
    .B1(_06398_),
    .Y(_06399_));
 sky130_fd_sc_hd__or2_1 _13711_ (.A(_06372_),
    .B(_06399_),
    .X(_06400_));
 sky130_fd_sc_hd__xnor2_1 _13712_ (.A(_06363_),
    .B(_06361_),
    .Y(_06401_));
 sky130_fd_sc_hd__xor2_2 _13713_ (.A(_06400_),
    .B(_06401_),
    .X(_06402_));
 sky130_fd_sc_hd__nor2_1 _13714_ (.A(_06383_),
    .B(_06397_),
    .Y(_06403_));
 sky130_fd_sc_hd__or2_1 _13715_ (.A(_06398_),
    .B(_06403_),
    .X(_06404_));
 sky130_fd_sc_hd__xnor2_2 _13716_ (.A(_06385_),
    .B(_06393_),
    .Y(_06405_));
 sky130_fd_sc_hd__and2_1 _13717_ (.A(_05641_),
    .B(_06304_),
    .X(_06406_));
 sky130_fd_sc_hd__clkbuf_2 _13718_ (.A(_06406_),
    .X(_06407_));
 sky130_fd_sc_hd__nand2_1 _13719_ (.A(_05738_),
    .B(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__xnor2_1 _13720_ (.A(_06327_),
    .B(_06378_),
    .Y(_06409_));
 sky130_fd_sc_hd__xor2_1 _13721_ (.A(_06408_),
    .B(_06409_),
    .X(_06410_));
 sky130_fd_sc_hd__and3_1 _13722_ (.A(_05567_),
    .B(_05748_),
    .C(_06320_),
    .X(_06411_));
 sky130_fd_sc_hd__or2_1 _13723_ (.A(_06266_),
    .B(_06331_),
    .X(_06412_));
 sky130_fd_sc_hd__xor2_1 _13724_ (.A(_06326_),
    .B(_06411_),
    .X(_06413_));
 sky130_fd_sc_hd__or2b_1 _13725_ (.A(_06412_),
    .B_N(_06413_),
    .X(_06414_));
 sky130_fd_sc_hd__a21boi_1 _13726_ (.A1(_06326_),
    .A2(_06411_),
    .B1_N(_06414_),
    .Y(_06415_));
 sky130_fd_sc_hd__or2b_1 _13727_ (.A(_06408_),
    .B_N(_06409_),
    .X(_06416_));
 sky130_fd_sc_hd__o21a_1 _13728_ (.A1(_06410_),
    .A2(_06415_),
    .B1(_06416_),
    .X(_06417_));
 sky130_fd_sc_hd__xnor2_2 _13729_ (.A(_06405_),
    .B(_06417_),
    .Y(_06418_));
 sky130_fd_sc_hd__o21bai_1 _13730_ (.A1(_05861_),
    .A2(_06389_),
    .B1_N(_06391_),
    .Y(_06419_));
 sky130_fd_sc_hd__nand2_1 _13731_ (.A(_06392_),
    .B(_06419_),
    .Y(_06420_));
 sky130_fd_sc_hd__nand2_1 _13732_ (.A(_06166_),
    .B(_06174_),
    .Y(_06421_));
 sky130_fd_sc_hd__nand2_2 _13733_ (.A(_06175_),
    .B(_06421_),
    .Y(_06422_));
 sky130_fd_sc_hd__clkbuf_4 _13734_ (.A(_06422_),
    .X(_06423_));
 sky130_fd_sc_hd__or2_1 _13735_ (.A(_05861_),
    .B(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__nor2_1 _13736_ (.A(_05767_),
    .B(_06343_),
    .Y(_06425_));
 sky130_fd_sc_hd__nor2_1 _13737_ (.A(_06317_),
    .B(_06388_),
    .Y(_06426_));
 sky130_fd_sc_hd__xnor2_1 _13738_ (.A(_06425_),
    .B(_06426_),
    .Y(_06427_));
 sky130_fd_sc_hd__nand2_1 _13739_ (.A(_06425_),
    .B(_06426_),
    .Y(_06428_));
 sky130_fd_sc_hd__o21a_1 _13740_ (.A1(_06424_),
    .A2(_06427_),
    .B1(_06428_),
    .X(_06429_));
 sky130_fd_sc_hd__o32ai_4 _13741_ (.A1(_06418_),
    .A2(_06420_),
    .A3(_06429_),
    .B1(_06417_),
    .B2(_06405_),
    .Y(_06430_));
 sky130_fd_sc_hd__and2_1 _13742_ (.A(_06374_),
    .B(_06394_),
    .X(_06431_));
 sky130_fd_sc_hd__or2_1 _13743_ (.A(_06395_),
    .B(_06431_),
    .X(_06432_));
 sky130_fd_sc_hd__nor2_1 _13744_ (.A(_06420_),
    .B(_06429_),
    .Y(_06433_));
 sky130_fd_sc_hd__xnor2_1 _13745_ (.A(_06418_),
    .B(_06433_),
    .Y(_06434_));
 sky130_fd_sc_hd__clkbuf_4 _13746_ (.A(_05638_),
    .X(_06435_));
 sky130_fd_sc_hd__and2_1 _13747_ (.A(_06376_),
    .B(_06379_),
    .X(_06436_));
 sky130_fd_sc_hd__or2_1 _13748_ (.A(_06380_),
    .B(_06436_),
    .X(_06437_));
 sky130_fd_sc_hd__o21ai_1 _13749_ (.A1(_06435_),
    .A2(_06306_),
    .B1(_06437_),
    .Y(_06438_));
 sky130_fd_sc_hd__xnor2_1 _13750_ (.A(_06410_),
    .B(_06415_),
    .Y(_06439_));
 sky130_fd_sc_hd__nand2_1 _13751_ (.A(_05738_),
    .B(_06305_),
    .Y(_06440_));
 sky130_fd_sc_hd__o21ai_1 _13752_ (.A1(_05740_),
    .A2(_06312_),
    .B1(_06440_),
    .Y(_06441_));
 sky130_fd_sc_hd__or2b_1 _13753_ (.A(_06439_),
    .B_N(_06441_),
    .X(_06442_));
 sky130_fd_sc_hd__xnor2_1 _13754_ (.A(_06438_),
    .B(_06442_),
    .Y(_06443_));
 sky130_fd_sc_hd__or2b_1 _13755_ (.A(_06442_),
    .B_N(_06438_),
    .X(_06444_));
 sky130_fd_sc_hd__a21boi_1 _13756_ (.A1(_06434_),
    .A2(_06443_),
    .B1_N(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__nor2_1 _13757_ (.A(_06432_),
    .B(_06445_),
    .Y(_06446_));
 sky130_fd_sc_hd__and2_1 _13758_ (.A(_06432_),
    .B(_06445_),
    .X(_06447_));
 sky130_fd_sc_hd__nor2_1 _13759_ (.A(_06446_),
    .B(_06447_),
    .Y(_06448_));
 sky130_fd_sc_hd__a21oi_1 _13760_ (.A1(_06430_),
    .A2(_06448_),
    .B1(_06446_),
    .Y(_06449_));
 sky130_fd_sc_hd__nor2_1 _13761_ (.A(_06404_),
    .B(_06449_),
    .Y(_06450_));
 sky130_fd_sc_hd__nand2_1 _13762_ (.A(_06372_),
    .B(_06399_),
    .Y(_06451_));
 sky130_fd_sc_hd__and2_1 _13763_ (.A(_06400_),
    .B(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__nand2_1 _13764_ (.A(_06450_),
    .B(_06452_),
    .Y(_06453_));
 sky130_fd_sc_hd__or2_1 _13765_ (.A(_06450_),
    .B(_06452_),
    .X(_06454_));
 sky130_fd_sc_hd__and2_1 _13766_ (.A(_06453_),
    .B(_06454_),
    .X(_06455_));
 sky130_fd_sc_hd__xnor2_1 _13767_ (.A(_06430_),
    .B(_06448_),
    .Y(_06456_));
 sky130_fd_sc_hd__xnor2_1 _13768_ (.A(_06434_),
    .B(_06443_),
    .Y(_06457_));
 sky130_fd_sc_hd__xor2_1 _13769_ (.A(_06441_),
    .B(_06439_),
    .X(_06458_));
 sky130_fd_sc_hd__xnor2_1 _13770_ (.A(_06412_),
    .B(_06413_),
    .Y(_06459_));
 sky130_fd_sc_hd__xor2_1 _13771_ (.A(_06408_),
    .B(_06459_),
    .X(_06460_));
 sky130_fd_sc_hd__nor2_1 _13772_ (.A(_06313_),
    .B(_06330_),
    .Y(_06461_));
 sky130_fd_sc_hd__nand3_1 _13773_ (.A(_06115_),
    .B(_06320_),
    .C(_06461_),
    .Y(_06462_));
 sky130_fd_sc_hd__nor2_1 _13774_ (.A(_06266_),
    .B(_06343_),
    .Y(_06463_));
 sky130_fd_sc_hd__a21o_1 _13775_ (.A1(_06115_),
    .A2(_06320_),
    .B1(_06461_),
    .X(_06464_));
 sky130_fd_sc_hd__nand3_1 _13776_ (.A(_06462_),
    .B(_06463_),
    .C(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__and2_1 _13777_ (.A(_06462_),
    .B(_06465_),
    .X(_06466_));
 sky130_fd_sc_hd__xor2_1 _13778_ (.A(_06460_),
    .B(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__xnor2_1 _13779_ (.A(_06440_),
    .B(_06407_),
    .Y(_06468_));
 sky130_fd_sc_hd__a211o_1 _13780_ (.A1(_05651_),
    .A2(_06311_),
    .B1(_06468_),
    .C1(_05434_),
    .X(_06469_));
 sky130_fd_sc_hd__buf_2 _13781_ (.A(_05660_),
    .X(_06470_));
 sky130_fd_sc_hd__a211o_1 _13782_ (.A1(_06260_),
    .A2(_06289_),
    .B1(_06303_),
    .C1(_06101_),
    .X(_06471_));
 sky130_fd_sc_hd__a211o_1 _13783_ (.A1(_06260_),
    .A2(_06289_),
    .B1(_06303_),
    .C1(_06470_),
    .X(_06472_));
 sky130_fd_sc_hd__a21boi_1 _13784_ (.A1(_05662_),
    .A2(_06471_),
    .B1_N(_06472_),
    .Y(_06473_));
 sky130_fd_sc_hd__a2bb2o_1 _13785_ (.A1_N(_06470_),
    .A2_N(_06471_),
    .B1(_06473_),
    .B2(_06468_),
    .X(_06474_));
 sky130_fd_sc_hd__or2_1 _13786_ (.A(_06469_),
    .B(_06474_),
    .X(_06475_));
 sky130_fd_sc_hd__nand2_1 _13787_ (.A(_06469_),
    .B(_06474_),
    .Y(_06476_));
 sky130_fd_sc_hd__a21boi_1 _13788_ (.A1(_06467_),
    .A2(_06475_),
    .B1_N(_06476_),
    .Y(_06477_));
 sky130_fd_sc_hd__xnor2_1 _13789_ (.A(_06424_),
    .B(_06427_),
    .Y(_06478_));
 sky130_fd_sc_hd__or2_1 _13790_ (.A(_05767_),
    .B(_06422_),
    .X(_06479_));
 sky130_fd_sc_hd__inv_2 _13791_ (.A(_06479_),
    .Y(_06480_));
 sky130_fd_sc_hd__nor2_1 _13792_ (.A(_06167_),
    .B(_06173_),
    .Y(_06481_));
 sky130_fd_sc_hd__nor2_1 _13793_ (.A(_06174_),
    .B(_06481_),
    .Y(_06482_));
 sky130_fd_sc_hd__buf_2 _13794_ (.A(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__or2_1 _13795_ (.A(_05861_),
    .B(_06483_),
    .X(_06484_));
 sky130_fd_sc_hd__o22a_1 _13796_ (.A1(_05767_),
    .A2(_06388_),
    .B1(_06422_),
    .B2(_06317_),
    .X(_06485_));
 sky130_fd_sc_hd__a21oi_1 _13797_ (.A1(_06426_),
    .A2(_06480_),
    .B1(_06485_),
    .Y(_06486_));
 sky130_fd_sc_hd__clkinv_2 _13798_ (.A(_06486_),
    .Y(_06487_));
 sky130_fd_sc_hd__o2bb2a_1 _13799_ (.A1_N(_06426_),
    .A2_N(_06480_),
    .B1(_06484_),
    .B2(_06487_),
    .X(_06488_));
 sky130_fd_sc_hd__or2_1 _13800_ (.A(_06478_),
    .B(_06488_),
    .X(_06489_));
 sky130_fd_sc_hd__and2_1 _13801_ (.A(_06420_),
    .B(_06429_),
    .X(_06490_));
 sky130_fd_sc_hd__or2_1 _13802_ (.A(_06433_),
    .B(_06490_),
    .X(_06491_));
 sky130_fd_sc_hd__or2b_1 _13803_ (.A(_06408_),
    .B_N(_06459_),
    .X(_06492_));
 sky130_fd_sc_hd__o21a_1 _13804_ (.A1(_06460_),
    .A2(_06466_),
    .B1(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__xor2_1 _13805_ (.A(_06491_),
    .B(_06493_),
    .X(_06494_));
 sky130_fd_sc_hd__xnor2_1 _13806_ (.A(_06489_),
    .B(_06494_),
    .Y(_06495_));
 sky130_fd_sc_hd__xor2_1 _13807_ (.A(_06458_),
    .B(_06477_),
    .X(_06496_));
 sky130_fd_sc_hd__nand2_1 _13808_ (.A(_06495_),
    .B(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__o21a_1 _13809_ (.A1(_06458_),
    .A2(_06477_),
    .B1(_06497_),
    .X(_06498_));
 sky130_fd_sc_hd__xnor2_1 _13810_ (.A(_06457_),
    .B(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__or2b_1 _13811_ (.A(_06489_),
    .B_N(_06494_),
    .X(_06500_));
 sky130_fd_sc_hd__o21ai_1 _13812_ (.A1(_06491_),
    .A2(_06493_),
    .B1(_06500_),
    .Y(_06501_));
 sky130_fd_sc_hd__or2b_1 _13813_ (.A(_06499_),
    .B_N(_06501_),
    .X(_06502_));
 sky130_fd_sc_hd__o21a_1 _13814_ (.A1(_06457_),
    .A2(_06498_),
    .B1(_06502_),
    .X(_06503_));
 sky130_fd_sc_hd__xor2_1 _13815_ (.A(_06456_),
    .B(_06503_),
    .X(_06504_));
 sky130_fd_sc_hd__xor2_1 _13816_ (.A(_06501_),
    .B(_06499_),
    .X(_06505_));
 sky130_fd_sc_hd__or2_1 _13817_ (.A(_06495_),
    .B(_06496_),
    .X(_06506_));
 sky130_fd_sc_hd__nand2_1 _13818_ (.A(_06497_),
    .B(_06506_),
    .Y(_06507_));
 sky130_fd_sc_hd__and2_1 _13819_ (.A(_06476_),
    .B(_06475_),
    .X(_06508_));
 sky130_fd_sc_hd__xnor2_1 _13820_ (.A(_06467_),
    .B(_06508_),
    .Y(_06509_));
 sky130_fd_sc_hd__nand2_2 _13821_ (.A(_05641_),
    .B(_06320_),
    .Y(_06510_));
 sky130_fd_sc_hd__a22o_1 _13822_ (.A1(_05641_),
    .A2(_06305_),
    .B1(_06321_),
    .B2(_05738_),
    .X(_06511_));
 sky130_fd_sc_hd__o21a_1 _13823_ (.A1(_06440_),
    .A2(_06510_),
    .B1(_06511_),
    .X(_06512_));
 sky130_fd_sc_hd__nand2_1 _13824_ (.A(_06471_),
    .B(_06472_),
    .Y(_06513_));
 sky130_fd_sc_hd__a21o_1 _13825_ (.A1(_05668_),
    .A2(_06311_),
    .B1(_06513_),
    .X(_06514_));
 sky130_fd_sc_hd__and2_1 _13826_ (.A(_05668_),
    .B(_06305_),
    .X(_06515_));
 sky130_fd_sc_hd__clkbuf_2 _13827_ (.A(_06515_),
    .X(_06516_));
 sky130_fd_sc_hd__xor2_1 _13828_ (.A(_06471_),
    .B(_06472_),
    .X(_06517_));
 sky130_fd_sc_hd__nand2_1 _13829_ (.A(_06516_),
    .B(_06517_),
    .Y(_06518_));
 sky130_fd_sc_hd__a21boi_1 _13830_ (.A1(_06512_),
    .A2(_06514_),
    .B1_N(_06518_),
    .Y(_06519_));
 sky130_fd_sc_hd__xor2_1 _13831_ (.A(_06468_),
    .B(_06473_),
    .X(_06520_));
 sky130_fd_sc_hd__or2b_1 _13832_ (.A(_06519_),
    .B_N(_06520_),
    .X(_06521_));
 sky130_fd_sc_hd__nor2_1 _13833_ (.A(_06440_),
    .B(_06510_),
    .Y(_06522_));
 sky130_fd_sc_hd__a21o_1 _13834_ (.A1(_06462_),
    .A2(_06464_),
    .B1(_06463_),
    .X(_06523_));
 sky130_fd_sc_hd__nand3_1 _13835_ (.A(_06465_),
    .B(_06522_),
    .C(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__a21o_1 _13836_ (.A1(_06465_),
    .A2(_06523_),
    .B1(_06522_),
    .X(_06525_));
 sky130_fd_sc_hd__or2_1 _13837_ (.A(_06310_),
    .B(_06342_),
    .X(_06526_));
 sky130_fd_sc_hd__or2_1 _13838_ (.A(_06310_),
    .B(_06330_),
    .X(_06527_));
 sky130_fd_sc_hd__nor2_1 _13839_ (.A(_06313_),
    .B(_06342_),
    .Y(_06528_));
 sky130_fd_sc_hd__xnor2_1 _13840_ (.A(_06527_),
    .B(_06528_),
    .Y(_06529_));
 sky130_fd_sc_hd__or3b_1 _13841_ (.A(_06266_),
    .B(_06389_),
    .C_N(_06529_),
    .X(_06530_));
 sky130_fd_sc_hd__o31ai_1 _13842_ (.A1(_06313_),
    .A2(_06331_),
    .A3(_06526_),
    .B1(_06530_),
    .Y(_06531_));
 sky130_fd_sc_hd__and3_1 _13843_ (.A(_06524_),
    .B(_06525_),
    .C(_06531_),
    .X(_06532_));
 sky130_fd_sc_hd__a21oi_1 _13844_ (.A1(_06524_),
    .A2(_06525_),
    .B1(_06531_),
    .Y(_06533_));
 sky130_fd_sc_hd__xor2_1 _13845_ (.A(_06520_),
    .B(_06519_),
    .X(_06534_));
 sky130_fd_sc_hd__or3_1 _13846_ (.A(_06532_),
    .B(_06533_),
    .C(_06534_),
    .X(_06535_));
 sky130_fd_sc_hd__nand2_1 _13847_ (.A(_06521_),
    .B(_06535_),
    .Y(_06536_));
 sky130_fd_sc_hd__and2b_1 _13848_ (.A_N(_06509_),
    .B(_06536_),
    .X(_06537_));
 sky130_fd_sc_hd__xor2_1 _13849_ (.A(_06484_),
    .B(_06486_),
    .X(_06538_));
 sky130_fd_sc_hd__or2_1 _13850_ (.A(_06317_),
    .B(_06483_),
    .X(_06539_));
 sky130_fd_sc_hd__or2_1 _13851_ (.A(_06168_),
    .B(_06172_),
    .X(_06540_));
 sky130_fd_sc_hd__nand2_1 _13852_ (.A(_06173_),
    .B(_06540_),
    .Y(_06541_));
 sky130_fd_sc_hd__buf_2 _13853_ (.A(_06541_),
    .X(_06542_));
 sky130_fd_sc_hd__or2_1 _13854_ (.A(_05861_),
    .B(_06542_),
    .X(_06543_));
 sky130_fd_sc_hd__xor2_1 _13855_ (.A(_06479_),
    .B(_06539_),
    .X(_06544_));
 sky130_fd_sc_hd__or2b_1 _13856_ (.A(_06543_),
    .B_N(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__o21a_1 _13857_ (.A1(_06479_),
    .A2(_06539_),
    .B1(_06545_),
    .X(_06546_));
 sky130_fd_sc_hd__nor2_1 _13858_ (.A(_06538_),
    .B(_06546_),
    .Y(_06547_));
 sky130_fd_sc_hd__a31o_1 _13859_ (.A1(_06465_),
    .A2(_06522_),
    .A3(_06523_),
    .B1(_06532_),
    .X(_06548_));
 sky130_fd_sc_hd__nand2_1 _13860_ (.A(_06478_),
    .B(_06488_),
    .Y(_06549_));
 sky130_fd_sc_hd__and2_1 _13861_ (.A(_06489_),
    .B(_06549_),
    .X(_06550_));
 sky130_fd_sc_hd__nor2_1 _13862_ (.A(_05434_),
    .B(_06550_),
    .Y(_06551_));
 sky130_fd_sc_hd__xnor2_1 _13863_ (.A(_06548_),
    .B(_06551_),
    .Y(_06552_));
 sky130_fd_sc_hd__xnor2_1 _13864_ (.A(_06547_),
    .B(_06552_),
    .Y(_06553_));
 sky130_fd_sc_hd__xnor2_1 _13865_ (.A(_06509_),
    .B(_06536_),
    .Y(_06554_));
 sky130_fd_sc_hd__and2b_1 _13866_ (.A_N(_06553_),
    .B(_06554_),
    .X(_06555_));
 sky130_fd_sc_hd__nor2_1 _13867_ (.A(_06537_),
    .B(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__xnor2_1 _13868_ (.A(_06507_),
    .B(_06556_),
    .Y(_06557_));
 sky130_fd_sc_hd__o21ai_1 _13869_ (.A1(_05434_),
    .A2(_06550_),
    .B1(_06548_),
    .Y(_06558_));
 sky130_fd_sc_hd__a21bo_1 _13870_ (.A1(_06547_),
    .A2(_06552_),
    .B1_N(_06558_),
    .X(_06559_));
 sky130_fd_sc_hd__or2b_1 _13871_ (.A(_06557_),
    .B_N(_06559_),
    .X(_06560_));
 sky130_fd_sc_hd__o21a_1 _13872_ (.A1(_06507_),
    .A2(_06556_),
    .B1(_06560_),
    .X(_06561_));
 sky130_fd_sc_hd__nor2_1 _13873_ (.A(_06505_),
    .B(_06561_),
    .Y(_06562_));
 sky130_fd_sc_hd__nand2_1 _13874_ (.A(_06504_),
    .B(_06562_),
    .Y(_06563_));
 sky130_fd_sc_hd__nor2_1 _13875_ (.A(_06456_),
    .B(_06503_),
    .Y(_06564_));
 sky130_fd_sc_hd__and2_1 _13876_ (.A(_06404_),
    .B(_06449_),
    .X(_06565_));
 sky130_fd_sc_hd__nor2_1 _13877_ (.A(_06450_),
    .B(_06565_),
    .Y(_06566_));
 sky130_fd_sc_hd__and2_1 _13878_ (.A(_06564_),
    .B(_06566_),
    .X(_06567_));
 sky130_fd_sc_hd__nor2_1 _13879_ (.A(_06564_),
    .B(_06566_),
    .Y(_06568_));
 sky130_fd_sc_hd__nor3_1 _13880_ (.A(_06563_),
    .B(_06567_),
    .C(_06568_),
    .Y(_06569_));
 sky130_fd_sc_hd__o21a_1 _13881_ (.A1(_06567_),
    .A2(_06568_),
    .B1(_06563_),
    .X(_06570_));
 sky130_fd_sc_hd__nor2_1 _13882_ (.A(_06569_),
    .B(_06570_),
    .Y(_06571_));
 sky130_fd_sc_hd__or2_1 _13883_ (.A(_06504_),
    .B(_06562_),
    .X(_06572_));
 sky130_fd_sc_hd__nand2_1 _13884_ (.A(_06563_),
    .B(_06572_),
    .Y(_06573_));
 sky130_fd_sc_hd__xor2_1 _13885_ (.A(_06505_),
    .B(_06561_),
    .X(_06574_));
 sky130_fd_sc_hd__xor2_1 _13886_ (.A(_06559_),
    .B(_06557_),
    .X(_06575_));
 sky130_fd_sc_hd__xor2_1 _13887_ (.A(_06553_),
    .B(_06554_),
    .X(_06576_));
 sky130_fd_sc_hd__xor2_1 _13888_ (.A(_06543_),
    .B(_06544_),
    .X(_06577_));
 sky130_fd_sc_hd__or2_1 _13889_ (.A(_05767_),
    .B(_06483_),
    .X(_06578_));
 sky130_fd_sc_hd__or2_1 _13890_ (.A(_06317_),
    .B(_06541_),
    .X(_06579_));
 sky130_fd_sc_hd__xnor2_1 _13891_ (.A(_06578_),
    .B(_06579_),
    .Y(_06580_));
 sky130_fd_sc_hd__or3_1 _13892_ (.A(_05861_),
    .B(_06172_),
    .C(_06580_),
    .X(_06581_));
 sky130_fd_sc_hd__o21a_1 _13893_ (.A1(_06578_),
    .A2(_06579_),
    .B1(_06581_),
    .X(_06582_));
 sky130_fd_sc_hd__or2_1 _13894_ (.A(_06577_),
    .B(_06582_),
    .X(_06583_));
 sky130_fd_sc_hd__and2_1 _13895_ (.A(_06538_),
    .B(_06546_),
    .X(_06584_));
 sky130_fd_sc_hd__or2_1 _13896_ (.A(_06547_),
    .B(_06584_),
    .X(_06585_));
 sky130_fd_sc_hd__or3_1 _13897_ (.A(_05434_),
    .B(_06137_),
    .C(_06305_),
    .X(_06586_));
 sky130_fd_sc_hd__nand2_1 _13898_ (.A(_06510_),
    .B(_06586_),
    .Y(_06587_));
 sky130_fd_sc_hd__nor2_1 _13899_ (.A(_06435_),
    .B(_06331_),
    .Y(_06588_));
 sky130_fd_sc_hd__nor2_1 _13900_ (.A(_06510_),
    .B(_06586_),
    .Y(_06589_));
 sky130_fd_sc_hd__a21o_1 _13901_ (.A1(_06587_),
    .A2(_06588_),
    .B1(_06589_),
    .X(_06590_));
 sky130_fd_sc_hd__a31o_1 _13902_ (.A1(_06230_),
    .A2(_06176_),
    .A3(_06387_),
    .B1(_06529_),
    .X(_06591_));
 sky130_fd_sc_hd__and2_1 _13903_ (.A(_06530_),
    .B(_06591_),
    .X(_06592_));
 sky130_fd_sc_hd__xnor2_1 _13904_ (.A(_06590_),
    .B(_06592_),
    .Y(_06593_));
 sky130_fd_sc_hd__nor2_1 _13905_ (.A(_06310_),
    .B(_06389_),
    .Y(_06594_));
 sky130_fd_sc_hd__nor2_1 _13906_ (.A(_06266_),
    .B(_06423_),
    .Y(_06595_));
 sky130_fd_sc_hd__nor2_1 _13907_ (.A(_06313_),
    .B(_06389_),
    .Y(_06596_));
 sky130_fd_sc_hd__xnor2_1 _13908_ (.A(_06526_),
    .B(_06596_),
    .Y(_06597_));
 sky130_fd_sc_hd__a22oi_2 _13909_ (.A1(_06528_),
    .A2(_06594_),
    .B1(_06595_),
    .B2(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__nand2_1 _13910_ (.A(_06590_),
    .B(_06592_),
    .Y(_06599_));
 sky130_fd_sc_hd__o21a_1 _13911_ (.A1(_06593_),
    .A2(_06598_),
    .B1(_06599_),
    .X(_06600_));
 sky130_fd_sc_hd__xor2_1 _13912_ (.A(_06585_),
    .B(_06600_),
    .X(_06601_));
 sky130_fd_sc_hd__xnor2_1 _13913_ (.A(_06583_),
    .B(_06601_),
    .Y(_06602_));
 sky130_fd_sc_hd__o21ai_1 _13914_ (.A1(_06532_),
    .A2(_06533_),
    .B1(_06534_),
    .Y(_06603_));
 sky130_fd_sc_hd__and2_1 _13915_ (.A(_06535_),
    .B(_06603_),
    .X(_06604_));
 sky130_fd_sc_hd__xor2_1 _13916_ (.A(_06593_),
    .B(_06598_),
    .X(_06605_));
 sky130_fd_sc_hd__nand2_1 _13917_ (.A(_06518_),
    .B(_06514_),
    .Y(_06606_));
 sky130_fd_sc_hd__xor2_1 _13918_ (.A(_06512_),
    .B(_06606_),
    .X(_06607_));
 sky130_fd_sc_hd__xnor2_1 _13919_ (.A(_06510_),
    .B(_06586_),
    .Y(_06608_));
 sky130_fd_sc_hd__xnor2_1 _13920_ (.A(_06608_),
    .B(_06588_),
    .Y(_06609_));
 sky130_fd_sc_hd__xnor2_1 _13921_ (.A(_06516_),
    .B(_06517_),
    .Y(_06610_));
 sky130_fd_sc_hd__a21bo_1 _13922_ (.A1(_05651_),
    .A2(_06320_),
    .B1_N(_06472_),
    .X(_06611_));
 sky130_fd_sc_hd__or3b_1 _13923_ (.A(_06471_),
    .B(_06470_),
    .C_N(_06320_),
    .X(_06612_));
 sky130_fd_sc_hd__a21bo_1 _13924_ (.A1(_06516_),
    .A2(_06611_),
    .B1_N(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__xnor2_1 _13925_ (.A(_06610_),
    .B(_06613_),
    .Y(_06614_));
 sky130_fd_sc_hd__and2b_1 _13926_ (.A_N(_06610_),
    .B(_06613_),
    .X(_06615_));
 sky130_fd_sc_hd__a21oi_1 _13927_ (.A1(_06609_),
    .A2(_06614_),
    .B1(_06615_),
    .Y(_06616_));
 sky130_fd_sc_hd__xor2_1 _13928_ (.A(_06607_),
    .B(_06616_),
    .X(_06617_));
 sky130_fd_sc_hd__nor2_1 _13929_ (.A(_06607_),
    .B(_06616_),
    .Y(_06618_));
 sky130_fd_sc_hd__a21oi_1 _13930_ (.A1(_06605_),
    .A2(_06617_),
    .B1(_06618_),
    .Y(_06619_));
 sky130_fd_sc_hd__xnor2_1 _13931_ (.A(_06604_),
    .B(_06619_),
    .Y(_06620_));
 sky130_fd_sc_hd__or2b_1 _13932_ (.A(_06619_),
    .B_N(_06604_),
    .X(_06621_));
 sky130_fd_sc_hd__a21boi_1 _13933_ (.A1(_06602_),
    .A2(_06620_),
    .B1_N(_06621_),
    .Y(_06622_));
 sky130_fd_sc_hd__xnor2_1 _13934_ (.A(_06576_),
    .B(_06622_),
    .Y(_06623_));
 sky130_fd_sc_hd__or2b_1 _13935_ (.A(_06583_),
    .B_N(_06601_),
    .X(_06624_));
 sky130_fd_sc_hd__o21ai_1 _13936_ (.A1(_06585_),
    .A2(_06600_),
    .B1(_06624_),
    .Y(_06625_));
 sky130_fd_sc_hd__or2b_1 _13937_ (.A(_06623_),
    .B_N(_06625_),
    .X(_06626_));
 sky130_fd_sc_hd__o21a_1 _13938_ (.A1(_06576_),
    .A2(_06622_),
    .B1(_06626_),
    .X(_06627_));
 sky130_fd_sc_hd__nor2_1 _13939_ (.A(_06575_),
    .B(_06627_),
    .Y(_06628_));
 sky130_fd_sc_hd__nand2_1 _13940_ (.A(_06574_),
    .B(_06628_),
    .Y(_06629_));
 sky130_fd_sc_hd__nand2_1 _13941_ (.A(_06573_),
    .B(_06629_),
    .Y(_06630_));
 sky130_fd_sc_hd__xnor2_1 _13942_ (.A(_06574_),
    .B(_06628_),
    .Y(_06631_));
 sky130_fd_sc_hd__xor2_1 _13943_ (.A(_06625_),
    .B(_06623_),
    .X(_06632_));
 sky130_fd_sc_hd__xnor2_1 _13944_ (.A(_06602_),
    .B(_06620_),
    .Y(_06633_));
 sky130_fd_sc_hd__buf_2 _13945_ (.A(_06172_),
    .X(_06634_));
 sky130_fd_sc_hd__or2_1 _13946_ (.A(_05767_),
    .B(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__nor2_1 _13947_ (.A(_06579_),
    .B(_06635_),
    .Y(_06636_));
 sky130_fd_sc_hd__o21ai_1 _13948_ (.A1(_05861_),
    .A2(_06634_),
    .B1(_06580_),
    .Y(_06637_));
 sky130_fd_sc_hd__and2_1 _13949_ (.A(_06581_),
    .B(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__nand2_1 _13950_ (.A(_06636_),
    .B(_06638_),
    .Y(_06639_));
 sky130_fd_sc_hd__nand2_1 _13951_ (.A(_06577_),
    .B(_06582_),
    .Y(_06640_));
 sky130_fd_sc_hd__nand2_1 _13952_ (.A(_06583_),
    .B(_06640_),
    .Y(_06641_));
 sky130_fd_sc_hd__nor2_1 _13953_ (.A(_06137_),
    .B(_06331_),
    .Y(_06642_));
 sky130_fd_sc_hd__nor2_1 _13954_ (.A(_05740_),
    .B(_06330_),
    .Y(_06643_));
 sky130_fd_sc_hd__a21o_1 _13955_ (.A1(_06028_),
    .A2(_06305_),
    .B1(_06643_),
    .X(_06644_));
 sky130_fd_sc_hd__nor2_1 _13956_ (.A(_06435_),
    .B(_06343_),
    .Y(_06645_));
 sky130_fd_sc_hd__a22o_1 _13957_ (.A1(_06407_),
    .A2(_06642_),
    .B1(_06644_),
    .B2(_06645_),
    .X(_06646_));
 sky130_fd_sc_hd__xor2_1 _13958_ (.A(_06595_),
    .B(_06597_),
    .X(_06647_));
 sky130_fd_sc_hd__xnor2_1 _13959_ (.A(_06646_),
    .B(_06647_),
    .Y(_06648_));
 sky130_fd_sc_hd__nor2_1 _13960_ (.A(_06310_),
    .B(_06423_),
    .Y(_06649_));
 sky130_fd_sc_hd__or2_1 _13961_ (.A(_06266_),
    .B(_06483_),
    .X(_06650_));
 sky130_fd_sc_hd__nor2_1 _13962_ (.A(_06313_),
    .B(_06422_),
    .Y(_06651_));
 sky130_fd_sc_hd__nor2_1 _13963_ (.A(_06594_),
    .B(_06651_),
    .Y(_06652_));
 sky130_fd_sc_hd__a21o_1 _13964_ (.A1(_06596_),
    .A2(_06649_),
    .B1(_06652_),
    .X(_06653_));
 sky130_fd_sc_hd__o2bb2a_1 _13965_ (.A1_N(_06596_),
    .A2_N(_06649_),
    .B1(_06650_),
    .B2(_06653_),
    .X(_06654_));
 sky130_fd_sc_hd__nor2_1 _13966_ (.A(_06648_),
    .B(_06654_),
    .Y(_06655_));
 sky130_fd_sc_hd__a21oi_1 _13967_ (.A1(_06646_),
    .A2(_06647_),
    .B1(_06655_),
    .Y(_06656_));
 sky130_fd_sc_hd__xor2_1 _13968_ (.A(_06641_),
    .B(_06656_),
    .X(_06657_));
 sky130_fd_sc_hd__xnor2_1 _13969_ (.A(_06639_),
    .B(_06657_),
    .Y(_06658_));
 sky130_fd_sc_hd__xnor2_1 _13970_ (.A(_06605_),
    .B(_06617_),
    .Y(_06659_));
 sky130_fd_sc_hd__and2_1 _13971_ (.A(_06648_),
    .B(_06654_),
    .X(_06660_));
 sky130_fd_sc_hd__nor2_1 _13972_ (.A(_06655_),
    .B(_06660_),
    .Y(_06661_));
 sky130_fd_sc_hd__xnor2_1 _13973_ (.A(_06609_),
    .B(_06614_),
    .Y(_06662_));
 sky130_fd_sc_hd__a21bo_1 _13974_ (.A1(_06407_),
    .A2(_06642_),
    .B1_N(_06644_),
    .X(_06663_));
 sky130_fd_sc_hd__xnor2_1 _13975_ (.A(_06663_),
    .B(_06645_),
    .Y(_06664_));
 sky130_fd_sc_hd__nand3_1 _13976_ (.A(_06516_),
    .B(_06612_),
    .C(_06611_),
    .Y(_06665_));
 sky130_fd_sc_hd__a21o_1 _13977_ (.A1(_06612_),
    .A2(_06611_),
    .B1(_06516_),
    .X(_06666_));
 sky130_fd_sc_hd__clkinv_2 _13978_ (.A(_06470_),
    .Y(_06667_));
 sky130_fd_sc_hd__a2bb2o_1 _13979_ (.A1_N(_06101_),
    .A2_N(_06331_),
    .B1(_06320_),
    .B2(_06667_),
    .X(_06668_));
 sky130_fd_sc_hd__nor2_1 _13980_ (.A(_06470_),
    .B(_06330_),
    .Y(_06669_));
 sky130_fd_sc_hd__nand3_1 _13981_ (.A(_05651_),
    .B(_06321_),
    .C(_06669_),
    .Y(_06670_));
 sky130_fd_sc_hd__a21bo_1 _13982_ (.A1(_06516_),
    .A2(_06668_),
    .B1_N(_06670_),
    .X(_06671_));
 sky130_fd_sc_hd__a21o_1 _13983_ (.A1(_06665_),
    .A2(_06666_),
    .B1(_06671_),
    .X(_06672_));
 sky130_fd_sc_hd__nand3_1 _13984_ (.A(_06665_),
    .B(_06666_),
    .C(_06671_),
    .Y(_06673_));
 sky130_fd_sc_hd__a21bo_1 _13985_ (.A1(_06664_),
    .A2(_06672_),
    .B1_N(_06673_),
    .X(_06674_));
 sky130_fd_sc_hd__xnor2_1 _13986_ (.A(_06662_),
    .B(_06674_),
    .Y(_06675_));
 sky130_fd_sc_hd__and2b_1 _13987_ (.A_N(_06662_),
    .B(_06674_),
    .X(_06676_));
 sky130_fd_sc_hd__a21oi_1 _13988_ (.A1(_06661_),
    .A2(_06675_),
    .B1(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__xor2_1 _13989_ (.A(_06659_),
    .B(_06677_),
    .X(_06678_));
 sky130_fd_sc_hd__nor2_1 _13990_ (.A(_06659_),
    .B(_06677_),
    .Y(_06679_));
 sky130_fd_sc_hd__a21oi_1 _13991_ (.A1(_06658_),
    .A2(_06678_),
    .B1(_06679_),
    .Y(_06680_));
 sky130_fd_sc_hd__xnor2_1 _13992_ (.A(_06633_),
    .B(_06680_),
    .Y(_06681_));
 sky130_fd_sc_hd__nor2_1 _13993_ (.A(_06641_),
    .B(_06656_),
    .Y(_06682_));
 sky130_fd_sc_hd__a31o_1 _13994_ (.A1(_06636_),
    .A2(_06638_),
    .A3(_06657_),
    .B1(_06682_),
    .X(_06683_));
 sky130_fd_sc_hd__or2b_1 _13995_ (.A(_06681_),
    .B_N(_06683_),
    .X(_06684_));
 sky130_fd_sc_hd__o21a_1 _13996_ (.A1(_06633_),
    .A2(_06680_),
    .B1(_06684_),
    .X(_06685_));
 sky130_fd_sc_hd__or2_1 _13997_ (.A(_06632_),
    .B(_06685_),
    .X(_06686_));
 sky130_fd_sc_hd__and2_1 _13998_ (.A(_06575_),
    .B(_06627_),
    .X(_06687_));
 sky130_fd_sc_hd__nor2_1 _13999_ (.A(_06628_),
    .B(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__and2b_1 _14000_ (.A_N(_06686_),
    .B(_06688_),
    .X(_06689_));
 sky130_fd_sc_hd__xnor2_1 _14001_ (.A(_06631_),
    .B(_06689_),
    .Y(_06690_));
 sky130_fd_sc_hd__nor2_1 _14002_ (.A(_06137_),
    .B(_06343_),
    .Y(_06691_));
 sky130_fd_sc_hd__a2bb2o_1 _14003_ (.A1_N(_05740_),
    .A2_N(_06343_),
    .B1(_06305_),
    .B2(_06028_),
    .X(_06692_));
 sky130_fd_sc_hd__nor2_1 _14004_ (.A(_05638_),
    .B(_06389_),
    .Y(_06693_));
 sky130_fd_sc_hd__a22o_1 _14005_ (.A1(_06407_),
    .A2(_06691_),
    .B1(_06692_),
    .B2(_06693_),
    .X(_06694_));
 sky130_fd_sc_hd__xor2_1 _14006_ (.A(_06650_),
    .B(_06653_),
    .X(_06695_));
 sky130_fd_sc_hd__nand2_1 _14007_ (.A(_06694_),
    .B(_06695_),
    .Y(_06696_));
 sky130_fd_sc_hd__xnor2_1 _14008_ (.A(_06694_),
    .B(_06695_),
    .Y(_06697_));
 sky130_fd_sc_hd__nor2_1 _14009_ (.A(_06310_),
    .B(_06483_),
    .Y(_06698_));
 sky130_fd_sc_hd__or2_1 _14010_ (.A(_06266_),
    .B(_06542_),
    .X(_06699_));
 sky130_fd_sc_hd__nor2_1 _14011_ (.A(_06313_),
    .B(_06483_),
    .Y(_06700_));
 sky130_fd_sc_hd__xnor2_1 _14012_ (.A(_06649_),
    .B(_06700_),
    .Y(_06701_));
 sky130_fd_sc_hd__o2bb2a_1 _14013_ (.A1_N(_06651_),
    .A2_N(_06698_),
    .B1(_06699_),
    .B2(_06701_),
    .X(_06702_));
 sky130_fd_sc_hd__or2_1 _14014_ (.A(_06697_),
    .B(_06702_),
    .X(_06703_));
 sky130_fd_sc_hd__or2_1 _14015_ (.A(_06636_),
    .B(_06638_),
    .X(_06704_));
 sky130_fd_sc_hd__nand2_1 _14016_ (.A(_06639_),
    .B(_06704_),
    .Y(_06705_));
 sky130_fd_sc_hd__a21oi_2 _14017_ (.A1(_06696_),
    .A2(_06703_),
    .B1(_06705_),
    .Y(_06706_));
 sky130_fd_sc_hd__xnor2_1 _14018_ (.A(_06658_),
    .B(_06678_),
    .Y(_06707_));
 sky130_fd_sc_hd__and3_1 _14019_ (.A(_06696_),
    .B(_06703_),
    .C(_06705_),
    .X(_06708_));
 sky130_fd_sc_hd__nor2_1 _14020_ (.A(_06706_),
    .B(_06708_),
    .Y(_06709_));
 sky130_fd_sc_hd__xnor2_1 _14021_ (.A(_06661_),
    .B(_06675_),
    .Y(_06710_));
 sky130_fd_sc_hd__nand2_1 _14022_ (.A(_06697_),
    .B(_06702_),
    .Y(_06711_));
 sky130_fd_sc_hd__and2_1 _14023_ (.A(_06703_),
    .B(_06711_),
    .X(_06712_));
 sky130_fd_sc_hd__nand3_1 _14024_ (.A(_06673_),
    .B(_06664_),
    .C(_06672_),
    .Y(_06713_));
 sky130_fd_sc_hd__a21o_1 _14025_ (.A1(_06673_),
    .A2(_06672_),
    .B1(_06664_),
    .X(_06714_));
 sky130_fd_sc_hd__a21bo_1 _14026_ (.A1(_06407_),
    .A2(_06691_),
    .B1_N(_06692_),
    .X(_06715_));
 sky130_fd_sc_hd__xnor2_1 _14027_ (.A(_06715_),
    .B(_06693_),
    .Y(_06716_));
 sky130_fd_sc_hd__nand3_1 _14028_ (.A(_06516_),
    .B(_06670_),
    .C(_06668_),
    .Y(_06717_));
 sky130_fd_sc_hd__a21o_1 _14029_ (.A1(_06670_),
    .A2(_06668_),
    .B1(_06516_),
    .X(_06718_));
 sky130_fd_sc_hd__nor2_1 _14030_ (.A(_06101_),
    .B(_06342_),
    .Y(_06719_));
 sky130_fd_sc_hd__xor2_1 _14031_ (.A(_06669_),
    .B(_06719_),
    .X(_06720_));
 sky130_fd_sc_hd__and2_1 _14032_ (.A(_06669_),
    .B(_06719_),
    .X(_06721_));
 sky130_fd_sc_hd__a31o_1 _14033_ (.A1(_05668_),
    .A2(_06321_),
    .A3(_06720_),
    .B1(_06721_),
    .X(_06722_));
 sky130_fd_sc_hd__a21o_1 _14034_ (.A1(_06717_),
    .A2(_06718_),
    .B1(_06722_),
    .X(_06723_));
 sky130_fd_sc_hd__nand3_1 _14035_ (.A(_06717_),
    .B(_06718_),
    .C(_06722_),
    .Y(_06724_));
 sky130_fd_sc_hd__a21bo_1 _14036_ (.A1(_06716_),
    .A2(_06723_),
    .B1_N(_06724_),
    .X(_06725_));
 sky130_fd_sc_hd__a21o_1 _14037_ (.A1(_06713_),
    .A2(_06714_),
    .B1(_06725_),
    .X(_06726_));
 sky130_fd_sc_hd__nand3_1 _14038_ (.A(_06713_),
    .B(_06714_),
    .C(_06725_),
    .Y(_06727_));
 sky130_fd_sc_hd__a21bo_1 _14039_ (.A1(_06712_),
    .A2(_06726_),
    .B1_N(_06727_),
    .X(_06728_));
 sky130_fd_sc_hd__xnor2_1 _14040_ (.A(_06710_),
    .B(_06728_),
    .Y(_06729_));
 sky130_fd_sc_hd__and2b_1 _14041_ (.A_N(_06710_),
    .B(_06728_),
    .X(_06730_));
 sky130_fd_sc_hd__a21oi_1 _14042_ (.A1(_06709_),
    .A2(_06729_),
    .B1(_06730_),
    .Y(_06731_));
 sky130_fd_sc_hd__xor2_2 _14043_ (.A(_06707_),
    .B(_06731_),
    .X(_06732_));
 sky130_fd_sc_hd__xnor2_2 _14044_ (.A(_06706_),
    .B(_06732_),
    .Y(_06733_));
 sky130_fd_sc_hd__and2_1 _14045_ (.A(_06028_),
    .B(_06305_),
    .X(_06734_));
 sky130_fd_sc_hd__nor2_1 _14046_ (.A(_05740_),
    .B(_06389_),
    .Y(_06735_));
 sky130_fd_sc_hd__xnor2_1 _14047_ (.A(_06734_),
    .B(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__nand2_1 _14048_ (.A(_06734_),
    .B(_06735_),
    .Y(_06737_));
 sky130_fd_sc_hd__o31ai_2 _14049_ (.A1(_06435_),
    .A2(_06423_),
    .A3(_06736_),
    .B1(_06737_),
    .Y(_06738_));
 sky130_fd_sc_hd__xor2_1 _14050_ (.A(_06699_),
    .B(_06701_),
    .X(_06739_));
 sky130_fd_sc_hd__nand2_1 _14051_ (.A(_06738_),
    .B(_06739_),
    .Y(_06740_));
 sky130_fd_sc_hd__xnor2_1 _14052_ (.A(_06738_),
    .B(_06739_),
    .Y(_06741_));
 sky130_fd_sc_hd__nor2_1 _14053_ (.A(_06313_),
    .B(_06542_),
    .Y(_06742_));
 sky130_fd_sc_hd__nor2_1 _14054_ (.A(_06310_),
    .B(_06542_),
    .Y(_06743_));
 sky130_fd_sc_hd__nor2_1 _14055_ (.A(_06698_),
    .B(_06742_),
    .Y(_06744_));
 sky130_fd_sc_hd__a21oi_1 _14056_ (.A1(_06700_),
    .A2(_06743_),
    .B1(_06744_),
    .Y(_06745_));
 sky130_fd_sc_hd__or3b_1 _14057_ (.A(_06266_),
    .B(_06172_),
    .C_N(_06745_),
    .X(_06746_));
 sky130_fd_sc_hd__a21boi_1 _14058_ (.A1(_06698_),
    .A2(_06742_),
    .B1_N(_06746_),
    .Y(_06747_));
 sky130_fd_sc_hd__or2_1 _14059_ (.A(_06741_),
    .B(_06747_),
    .X(_06748_));
 sky130_fd_sc_hd__o22a_1 _14060_ (.A1(_06317_),
    .A2(_06634_),
    .B1(_06542_),
    .B2(_05767_),
    .X(_06749_));
 sky130_fd_sc_hd__or2_1 _14061_ (.A(_06636_),
    .B(_06749_),
    .X(_06750_));
 sky130_fd_sc_hd__a21oi_2 _14062_ (.A1(_06740_),
    .A2(_06748_),
    .B1(_06750_),
    .Y(_06751_));
 sky130_fd_sc_hd__xnor2_1 _14063_ (.A(_06709_),
    .B(_06729_),
    .Y(_06752_));
 sky130_fd_sc_hd__and3_1 _14064_ (.A(_06740_),
    .B(_06748_),
    .C(_06750_),
    .X(_06753_));
 sky130_fd_sc_hd__nor2_1 _14065_ (.A(_06751_),
    .B(_06753_),
    .Y(_06754_));
 sky130_fd_sc_hd__nand3_1 _14066_ (.A(_06727_),
    .B(_06712_),
    .C(_06726_),
    .Y(_06755_));
 sky130_fd_sc_hd__a21o_1 _14067_ (.A1(_06727_),
    .A2(_06726_),
    .B1(_06712_),
    .X(_06756_));
 sky130_fd_sc_hd__xor2_1 _14068_ (.A(_06741_),
    .B(_06747_),
    .X(_06757_));
 sky130_fd_sc_hd__nand3_1 _14069_ (.A(_06724_),
    .B(_06716_),
    .C(_06723_),
    .Y(_06758_));
 sky130_fd_sc_hd__a21o_1 _14070_ (.A1(_06724_),
    .A2(_06723_),
    .B1(_06716_),
    .X(_06759_));
 sky130_fd_sc_hd__nor2_1 _14071_ (.A(_06435_),
    .B(_06423_),
    .Y(_06760_));
 sky130_fd_sc_hd__xnor2_1 _14072_ (.A(_06736_),
    .B(_06760_),
    .Y(_06761_));
 sky130_fd_sc_hd__nand2_1 _14073_ (.A(_05668_),
    .B(_06321_),
    .Y(_06762_));
 sky130_fd_sc_hd__xnor2_1 _14074_ (.A(_06762_),
    .B(_06720_),
    .Y(_06763_));
 sky130_fd_sc_hd__nor2_1 _14075_ (.A(_06470_),
    .B(_06388_),
    .Y(_06764_));
 sky130_fd_sc_hd__nor2_1 _14076_ (.A(_05959_),
    .B(_06331_),
    .Y(_06765_));
 sky130_fd_sc_hd__or2_1 _14077_ (.A(_06470_),
    .B(_06342_),
    .X(_06766_));
 sky130_fd_sc_hd__nor2_1 _14078_ (.A(_06101_),
    .B(_06389_),
    .Y(_06767_));
 sky130_fd_sc_hd__xnor2_1 _14079_ (.A(_06766_),
    .B(_06767_),
    .Y(_06768_));
 sky130_fd_sc_hd__a22o_1 _14080_ (.A1(_06719_),
    .A2(_06764_),
    .B1(_06765_),
    .B2(_06768_),
    .X(_06769_));
 sky130_fd_sc_hd__xor2_1 _14081_ (.A(_06763_),
    .B(_06769_),
    .X(_06770_));
 sky130_fd_sc_hd__and2_1 _14082_ (.A(_06763_),
    .B(_06769_),
    .X(_06771_));
 sky130_fd_sc_hd__a21o_1 _14083_ (.A1(_06761_),
    .A2(_06770_),
    .B1(_06771_),
    .X(_06772_));
 sky130_fd_sc_hd__a21o_1 _14084_ (.A1(_06758_),
    .A2(_06759_),
    .B1(_06772_),
    .X(_06773_));
 sky130_fd_sc_hd__nand3_1 _14085_ (.A(_06758_),
    .B(_06759_),
    .C(_06772_),
    .Y(_06774_));
 sky130_fd_sc_hd__a21bo_1 _14086_ (.A1(_06757_),
    .A2(_06773_),
    .B1_N(_06774_),
    .X(_06775_));
 sky130_fd_sc_hd__a21o_1 _14087_ (.A1(_06755_),
    .A2(_06756_),
    .B1(_06775_),
    .X(_06776_));
 sky130_fd_sc_hd__nand3_1 _14088_ (.A(_06755_),
    .B(_06756_),
    .C(_06775_),
    .Y(_06777_));
 sky130_fd_sc_hd__a21bo_1 _14089_ (.A1(_06754_),
    .A2(_06776_),
    .B1_N(_06777_),
    .X(_06778_));
 sky130_fd_sc_hd__xnor2_1 _14090_ (.A(_06752_),
    .B(_06778_),
    .Y(_06779_));
 sky130_fd_sc_hd__and2b_1 _14091_ (.A_N(_06752_),
    .B(_06778_),
    .X(_06780_));
 sky130_fd_sc_hd__a21oi_2 _14092_ (.A1(_06751_),
    .A2(_06779_),
    .B1(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__nor2_1 _14093_ (.A(_06733_),
    .B(_06781_),
    .Y(_06782_));
 sky130_fd_sc_hd__or2_1 _14094_ (.A(_06707_),
    .B(_06731_),
    .X(_06783_));
 sky130_fd_sc_hd__nand2_1 _14095_ (.A(_06706_),
    .B(_06732_),
    .Y(_06784_));
 sky130_fd_sc_hd__xor2_1 _14096_ (.A(_06683_),
    .B(_06681_),
    .X(_06785_));
 sky130_fd_sc_hd__a21oi_1 _14097_ (.A1(_06783_),
    .A2(_06784_),
    .B1(_06785_),
    .Y(_06786_));
 sky130_fd_sc_hd__and3_1 _14098_ (.A(_06785_),
    .B(_06783_),
    .C(_06784_),
    .X(_06787_));
 sky130_fd_sc_hd__nor2_1 _14099_ (.A(_06786_),
    .B(_06787_),
    .Y(_06788_));
 sky130_fd_sc_hd__and2_1 _14100_ (.A(_06782_),
    .B(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__xor2_1 _14101_ (.A(_06632_),
    .B(_06685_),
    .X(_06790_));
 sky130_fd_sc_hd__and2_1 _14102_ (.A(_06786_),
    .B(_06790_),
    .X(_06791_));
 sky130_fd_sc_hd__nor2_1 _14103_ (.A(_06786_),
    .B(_06790_),
    .Y(_06792_));
 sky130_fd_sc_hd__nor2_1 _14104_ (.A(_06791_),
    .B(_06792_),
    .Y(_06793_));
 sky130_fd_sc_hd__or2_1 _14105_ (.A(_06789_),
    .B(_06793_),
    .X(_06794_));
 sky130_fd_sc_hd__xor2_2 _14106_ (.A(_06733_),
    .B(_06781_),
    .X(_06795_));
 sky130_fd_sc_hd__nand3_1 _14107_ (.A(_06777_),
    .B(_06754_),
    .C(_06776_),
    .Y(_06796_));
 sky130_fd_sc_hd__a21o_1 _14108_ (.A1(_06777_),
    .A2(_06776_),
    .B1(_06754_),
    .X(_06797_));
 sky130_fd_sc_hd__and2_1 _14109_ (.A(_05641_),
    .B(_06321_),
    .X(_06798_));
 sky130_fd_sc_hd__nor2_1 _14110_ (.A(_06137_),
    .B(_06423_),
    .Y(_06799_));
 sky130_fd_sc_hd__a2bb2o_1 _14111_ (.A1_N(_05740_),
    .A2_N(_06423_),
    .B1(_06321_),
    .B2(_06028_),
    .X(_06800_));
 sky130_fd_sc_hd__nor2_1 _14112_ (.A(_06435_),
    .B(_06483_),
    .Y(_06801_));
 sky130_fd_sc_hd__a22o_1 _14113_ (.A1(_06798_),
    .A2(_06799_),
    .B1(_06800_),
    .B2(_06801_),
    .X(_06802_));
 sky130_fd_sc_hd__o21bai_1 _14114_ (.A1(_06266_),
    .A2(_06634_),
    .B1_N(_06745_),
    .Y(_06803_));
 sky130_fd_sc_hd__nor2_1 _14115_ (.A(_06313_),
    .B(_06634_),
    .Y(_06804_));
 sky130_fd_sc_hd__nand2_1 _14116_ (.A(_06746_),
    .B(_06803_),
    .Y(_06805_));
 sky130_fd_sc_hd__xnor2_1 _14117_ (.A(_06802_),
    .B(_06805_),
    .Y(_06806_));
 sky130_fd_sc_hd__and3_1 _14118_ (.A(_06743_),
    .B(_06804_),
    .C(_06806_),
    .X(_06807_));
 sky130_fd_sc_hd__a31oi_1 _14119_ (.A1(_06746_),
    .A2(_06802_),
    .A3(_06803_),
    .B1(_06807_),
    .Y(_06808_));
 sky130_fd_sc_hd__nor2_1 _14120_ (.A(_06635_),
    .B(_06808_),
    .Y(_06809_));
 sky130_fd_sc_hd__and2_1 _14121_ (.A(_06635_),
    .B(_06808_),
    .X(_06810_));
 sky130_fd_sc_hd__nor2_1 _14122_ (.A(_06809_),
    .B(_06810_),
    .Y(_06811_));
 sky130_fd_sc_hd__nand3_1 _14123_ (.A(_06774_),
    .B(_06757_),
    .C(_06773_),
    .Y(_06812_));
 sky130_fd_sc_hd__a21o_1 _14124_ (.A1(_06774_),
    .A2(_06773_),
    .B1(_06757_),
    .X(_06813_));
 sky130_fd_sc_hd__xnor2_1 _14125_ (.A(_06761_),
    .B(_06770_),
    .Y(_06814_));
 sky130_fd_sc_hd__o31a_1 _14126_ (.A1(_06137_),
    .A2(_06423_),
    .A3(_06510_),
    .B1(_06800_),
    .X(_06815_));
 sky130_fd_sc_hd__xor2_1 _14127_ (.A(_06815_),
    .B(_06801_),
    .X(_06816_));
 sky130_fd_sc_hd__xnor2_1 _14128_ (.A(_06765_),
    .B(_06768_),
    .Y(_06817_));
 sky130_fd_sc_hd__nor2_1 _14129_ (.A(_06101_),
    .B(_06422_),
    .Y(_06818_));
 sky130_fd_sc_hd__xor2_1 _14130_ (.A(_06764_),
    .B(_06818_),
    .X(_06819_));
 sky130_fd_sc_hd__or3b_1 _14131_ (.A(_05959_),
    .B(_06343_),
    .C_N(_06819_),
    .X(_06820_));
 sky130_fd_sc_hd__a21bo_1 _14132_ (.A1(_06764_),
    .A2(_06818_),
    .B1_N(_06820_),
    .X(_06821_));
 sky130_fd_sc_hd__xnor2_1 _14133_ (.A(_06817_),
    .B(_06821_),
    .Y(_06822_));
 sky130_fd_sc_hd__and2b_1 _14134_ (.A_N(_06817_),
    .B(_06821_),
    .X(_06823_));
 sky130_fd_sc_hd__a21oi_1 _14135_ (.A1(_06816_),
    .A2(_06822_),
    .B1(_06823_),
    .Y(_06824_));
 sky130_fd_sc_hd__nor2_1 _14136_ (.A(_06814_),
    .B(_06824_),
    .Y(_06825_));
 sky130_fd_sc_hd__nor2_1 _14137_ (.A(_06310_),
    .B(_06634_),
    .Y(_06826_));
 sky130_fd_sc_hd__nand2_1 _14138_ (.A(_06742_),
    .B(_06826_),
    .Y(_06827_));
 sky130_fd_sc_hd__xor2_1 _14139_ (.A(_06827_),
    .B(_06806_),
    .X(_06828_));
 sky130_fd_sc_hd__inv_2 _14140_ (.A(_06828_),
    .Y(_06829_));
 sky130_fd_sc_hd__xor2_1 _14141_ (.A(_06814_),
    .B(_06824_),
    .X(_06830_));
 sky130_fd_sc_hd__and2_1 _14142_ (.A(_06829_),
    .B(_06830_),
    .X(_06831_));
 sky130_fd_sc_hd__a211o_1 _14143_ (.A1(_06812_),
    .A2(_06813_),
    .B1(_06825_),
    .C1(_06831_),
    .X(_06832_));
 sky130_fd_sc_hd__o211a_1 _14144_ (.A1(_06825_),
    .A2(_06831_),
    .B1(_06812_),
    .C1(_06813_),
    .X(_06833_));
 sky130_fd_sc_hd__a21o_1 _14145_ (.A1(_06811_),
    .A2(_06832_),
    .B1(_06833_),
    .X(_06834_));
 sky130_fd_sc_hd__nand3_1 _14146_ (.A(_06796_),
    .B(_06797_),
    .C(_06834_),
    .Y(_06835_));
 sky130_fd_sc_hd__inv_2 _14147_ (.A(_06835_),
    .Y(_06836_));
 sky130_fd_sc_hd__a21o_1 _14148_ (.A1(_06796_),
    .A2(_06797_),
    .B1(_06834_),
    .X(_06837_));
 sky130_fd_sc_hd__and3_1 _14149_ (.A(_06809_),
    .B(_06835_),
    .C(_06837_),
    .X(_06838_));
 sky130_fd_sc_hd__xnor2_1 _14150_ (.A(_06751_),
    .B(_06779_),
    .Y(_06839_));
 sky130_fd_sc_hd__o21ba_1 _14151_ (.A1(_06836_),
    .A2(_06838_),
    .B1_N(_06839_),
    .X(_06840_));
 sky130_fd_sc_hd__and2_1 _14152_ (.A(_06795_),
    .B(_06840_),
    .X(_06841_));
 sky130_fd_sc_hd__or2b_1 _14153_ (.A(_06833_),
    .B_N(_06832_),
    .X(_06842_));
 sky130_fd_sc_hd__xor2_1 _14154_ (.A(_06811_),
    .B(_06842_),
    .X(_06843_));
 sky130_fd_sc_hd__nor2_1 _14155_ (.A(_06137_),
    .B(_06483_),
    .Y(_06844_));
 sky130_fd_sc_hd__nand2_1 _14156_ (.A(_06643_),
    .B(_06844_),
    .Y(_06845_));
 sky130_fd_sc_hd__nor2_1 _14157_ (.A(_05740_),
    .B(_06483_),
    .Y(_06846_));
 sky130_fd_sc_hd__xnor2_1 _14158_ (.A(_06642_),
    .B(_06846_),
    .Y(_06847_));
 sky130_fd_sc_hd__or3_1 _14159_ (.A(_06435_),
    .B(_06542_),
    .C(_06847_),
    .X(_06848_));
 sky130_fd_sc_hd__or2_1 _14160_ (.A(_06743_),
    .B(_06804_),
    .X(_06849_));
 sky130_fd_sc_hd__nand2_1 _14161_ (.A(_06827_),
    .B(_06849_),
    .Y(_06850_));
 sky130_fd_sc_hd__a21o_1 _14162_ (.A1(_06845_),
    .A2(_06848_),
    .B1(_06850_),
    .X(_06851_));
 sky130_fd_sc_hd__nor2_1 _14163_ (.A(_06829_),
    .B(_06830_),
    .Y(_06852_));
 sky130_fd_sc_hd__or2_1 _14164_ (.A(_06831_),
    .B(_06852_),
    .X(_06853_));
 sky130_fd_sc_hd__nand3_1 _14165_ (.A(_06845_),
    .B(_06848_),
    .C(_06850_),
    .Y(_06854_));
 sky130_fd_sc_hd__and2_1 _14166_ (.A(_06851_),
    .B(_06854_),
    .X(_06855_));
 sky130_fd_sc_hd__a31o_1 _14167_ (.A1(_05668_),
    .A2(_06222_),
    .A3(_06341_),
    .B1(_06819_),
    .X(_06856_));
 sky130_fd_sc_hd__nand2_1 _14168_ (.A(_06820_),
    .B(_06856_),
    .Y(_06857_));
 sky130_fd_sc_hd__or2_1 _14169_ (.A(_05660_),
    .B(_06482_),
    .X(_06858_));
 sky130_fd_sc_hd__or2_1 _14170_ (.A(_06470_),
    .B(_06422_),
    .X(_06859_));
 sky130_fd_sc_hd__nor2_1 _14171_ (.A(_06101_),
    .B(_06482_),
    .Y(_06860_));
 sky130_fd_sc_hd__xnor2_1 _14172_ (.A(_06859_),
    .B(_06860_),
    .Y(_06861_));
 sky130_fd_sc_hd__or3b_1 _14173_ (.A(_05959_),
    .B(_06389_),
    .C_N(_06861_),
    .X(_06862_));
 sky130_fd_sc_hd__o31a_1 _14174_ (.A1(_06101_),
    .A2(_06423_),
    .A3(_06858_),
    .B1(_06862_),
    .X(_06863_));
 sky130_fd_sc_hd__o21ai_1 _14175_ (.A1(_06435_),
    .A2(_06542_),
    .B1(_06847_),
    .Y(_06864_));
 sky130_fd_sc_hd__nand2_1 _14176_ (.A(_06848_),
    .B(_06864_),
    .Y(_06865_));
 sky130_fd_sc_hd__xor2_1 _14177_ (.A(_06857_),
    .B(_06863_),
    .X(_06866_));
 sky130_fd_sc_hd__or2b_1 _14178_ (.A(_06865_),
    .B_N(_06866_),
    .X(_06867_));
 sky130_fd_sc_hd__o21a_1 _14179_ (.A1(_06857_),
    .A2(_06863_),
    .B1(_06867_),
    .X(_06868_));
 sky130_fd_sc_hd__xor2_1 _14180_ (.A(_06816_),
    .B(_06822_),
    .X(_06869_));
 sky130_fd_sc_hd__and2b_1 _14181_ (.A_N(_06868_),
    .B(_06869_),
    .X(_06870_));
 sky130_fd_sc_hd__and2b_1 _14182_ (.A_N(_06869_),
    .B(_06868_),
    .X(_06871_));
 sky130_fd_sc_hd__nor2_1 _14183_ (.A(_06870_),
    .B(_06871_),
    .Y(_06872_));
 sky130_fd_sc_hd__a21oi_1 _14184_ (.A1(_06855_),
    .A2(_06872_),
    .B1(_06870_),
    .Y(_06873_));
 sky130_fd_sc_hd__and2_1 _14185_ (.A(_06853_),
    .B(_06873_),
    .X(_06874_));
 sky130_fd_sc_hd__nor2_1 _14186_ (.A(_06853_),
    .B(_06873_),
    .Y(_06875_));
 sky130_fd_sc_hd__o21ba_1 _14187_ (.A1(_06851_),
    .A2(_06874_),
    .B1_N(_06875_),
    .X(_06876_));
 sky130_fd_sc_hd__nor2_1 _14188_ (.A(_06843_),
    .B(_06876_),
    .Y(_06877_));
 sky130_fd_sc_hd__a21oi_1 _14189_ (.A1(_06835_),
    .A2(_06837_),
    .B1(_06809_),
    .Y(_06878_));
 sky130_fd_sc_hd__a211oi_1 _14190_ (.A1(_06839_),
    .A2(_06835_),
    .B1(_06838_),
    .C1(_06878_),
    .Y(_06879_));
 sky130_fd_sc_hd__nand2_1 _14191_ (.A(_06843_),
    .B(_06876_),
    .Y(_06880_));
 sky130_fd_sc_hd__or2_1 _14192_ (.A(_05740_),
    .B(_06542_),
    .X(_06881_));
 sky130_fd_sc_hd__xor2_1 _14193_ (.A(_06691_),
    .B(_06881_),
    .X(_06882_));
 sky130_fd_sc_hd__or3_1 _14194_ (.A(_06137_),
    .B(_06343_),
    .C(_06881_),
    .X(_06883_));
 sky130_fd_sc_hd__o31a_1 _14195_ (.A1(_06435_),
    .A2(_06634_),
    .A3(_06882_),
    .B1(_06883_),
    .X(_06884_));
 sky130_fd_sc_hd__or3_1 _14196_ (.A(_06310_),
    .B(_06634_),
    .C(_06884_),
    .X(_06885_));
 sky130_fd_sc_hd__xnor2_1 _14197_ (.A(_06855_),
    .B(_06872_),
    .Y(_06886_));
 sky130_fd_sc_hd__xor2_1 _14198_ (.A(_06865_),
    .B(_06866_),
    .X(_06887_));
 sky130_fd_sc_hd__a31o_1 _14199_ (.A1(_05668_),
    .A2(_06176_),
    .A3(_06387_),
    .B1(_06861_),
    .X(_06888_));
 sky130_fd_sc_hd__or2_1 _14200_ (.A(_06101_),
    .B(_06541_),
    .X(_06889_));
 sky130_fd_sc_hd__xor2_1 _14201_ (.A(_06858_),
    .B(_06889_),
    .X(_06890_));
 sky130_fd_sc_hd__or3b_1 _14202_ (.A(_05959_),
    .B(_06423_),
    .C_N(_06890_),
    .X(_06891_));
 sky130_fd_sc_hd__o21ai_1 _14203_ (.A1(_06858_),
    .A2(_06889_),
    .B1(_06891_),
    .Y(_06892_));
 sky130_fd_sc_hd__nor2_1 _14204_ (.A(_06435_),
    .B(_06634_),
    .Y(_06893_));
 sky130_fd_sc_hd__xnor2_1 _14205_ (.A(_06882_),
    .B(_06893_),
    .Y(_06894_));
 sky130_fd_sc_hd__nand2_1 _14206_ (.A(_06862_),
    .B(_06888_),
    .Y(_06895_));
 sky130_fd_sc_hd__xnor2_1 _14207_ (.A(_06895_),
    .B(_06892_),
    .Y(_06896_));
 sky130_fd_sc_hd__a32o_1 _14208_ (.A1(_06862_),
    .A2(_06888_),
    .A3(_06892_),
    .B1(_06894_),
    .B2(_06896_),
    .X(_06897_));
 sky130_fd_sc_hd__or2b_1 _14209_ (.A(_06887_),
    .B_N(_06897_),
    .X(_06898_));
 sky130_fd_sc_hd__xnor2_1 _14210_ (.A(_06826_),
    .B(_06884_),
    .Y(_06899_));
 sky130_fd_sc_hd__xnor2_1 _14211_ (.A(_06887_),
    .B(_06897_),
    .Y(_06900_));
 sky130_fd_sc_hd__nand2_1 _14212_ (.A(_06899_),
    .B(_06900_),
    .Y(_06901_));
 sky130_fd_sc_hd__and2_1 _14213_ (.A(_06898_),
    .B(_06901_),
    .X(_06902_));
 sky130_fd_sc_hd__nor2_1 _14214_ (.A(_06886_),
    .B(_06902_),
    .Y(_06903_));
 sky130_fd_sc_hd__and2_1 _14215_ (.A(_06886_),
    .B(_06902_),
    .X(_06904_));
 sky130_fd_sc_hd__or2_1 _14216_ (.A(_06903_),
    .B(_06904_),
    .X(_06905_));
 sky130_fd_sc_hd__nand2_1 _14217_ (.A(_06885_),
    .B(_06905_),
    .Y(_06906_));
 sky130_fd_sc_hd__or2_1 _14218_ (.A(_06899_),
    .B(_06900_),
    .X(_06907_));
 sky130_fd_sc_hd__nand2_1 _14219_ (.A(_06901_),
    .B(_06907_),
    .Y(_06908_));
 sky130_fd_sc_hd__nand2_1 _14220_ (.A(_06894_),
    .B(_06896_),
    .Y(_06909_));
 sky130_fd_sc_hd__or2_1 _14221_ (.A(_06894_),
    .B(_06896_),
    .X(_06910_));
 sky130_fd_sc_hd__nand2_1 _14222_ (.A(_06909_),
    .B(_06910_),
    .Y(_06911_));
 sky130_fd_sc_hd__a31o_1 _14223_ (.A1(_05668_),
    .A2(_06175_),
    .A3(_06421_),
    .B1(_06890_),
    .X(_06912_));
 sky130_fd_sc_hd__nand2_1 _14224_ (.A(_06891_),
    .B(_06912_),
    .Y(_06913_));
 sky130_fd_sc_hd__or2_1 _14225_ (.A(_06470_),
    .B(_06172_),
    .X(_06914_));
 sky130_fd_sc_hd__nor2_1 _14226_ (.A(_05959_),
    .B(_06483_),
    .Y(_06915_));
 sky130_fd_sc_hd__o22a_1 _14227_ (.A1(_06101_),
    .A2(_06172_),
    .B1(_06542_),
    .B2(_06470_),
    .X(_06916_));
 sky130_fd_sc_hd__o21ba_1 _14228_ (.A1(_06889_),
    .A2(_06914_),
    .B1_N(_06916_),
    .X(_06917_));
 sky130_fd_sc_hd__a2bb2o_1 _14229_ (.A1_N(_06889_),
    .A2_N(_06914_),
    .B1(_06915_),
    .B2(_06917_),
    .X(_06918_));
 sky130_fd_sc_hd__inv_2 _14230_ (.A(_06918_),
    .Y(_06919_));
 sky130_fd_sc_hd__nor2_1 _14231_ (.A(_06137_),
    .B(_06172_),
    .Y(_06920_));
 sky130_fd_sc_hd__and2_1 _14232_ (.A(_06735_),
    .B(_06920_),
    .X(_06921_));
 sky130_fd_sc_hd__o22a_1 _14233_ (.A1(_05740_),
    .A2(_06634_),
    .B1(_06389_),
    .B2(_06137_),
    .X(_06922_));
 sky130_fd_sc_hd__nor2_1 _14234_ (.A(_06921_),
    .B(_06922_),
    .Y(_06923_));
 sky130_fd_sc_hd__xnor2_1 _14235_ (.A(_06913_),
    .B(_06918_),
    .Y(_06924_));
 sky130_fd_sc_hd__nand2_1 _14236_ (.A(_06923_),
    .B(_06924_),
    .Y(_06925_));
 sky130_fd_sc_hd__o21a_1 _14237_ (.A1(_06913_),
    .A2(_06919_),
    .B1(_06925_),
    .X(_06926_));
 sky130_fd_sc_hd__or2_1 _14238_ (.A(_06911_),
    .B(_06926_),
    .X(_06927_));
 sky130_fd_sc_hd__nand2_1 _14239_ (.A(_06911_),
    .B(_06926_),
    .Y(_06928_));
 sky130_fd_sc_hd__and2_1 _14240_ (.A(_06927_),
    .B(_06928_),
    .X(_06929_));
 sky130_fd_sc_hd__nand2_1 _14241_ (.A(_06921_),
    .B(_06929_),
    .Y(_06930_));
 sky130_fd_sc_hd__nand3_1 _14242_ (.A(_06908_),
    .B(_06927_),
    .C(_06930_),
    .Y(_06931_));
 sky130_fd_sc_hd__or2_1 _14243_ (.A(_06923_),
    .B(_06924_),
    .X(_06932_));
 sky130_fd_sc_hd__nand2_1 _14244_ (.A(_06925_),
    .B(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__or2_1 _14245_ (.A(_05959_),
    .B(_06542_),
    .X(_06934_));
 sky130_fd_sc_hd__or2_1 _14246_ (.A(_06914_),
    .B(_06934_),
    .X(_06935_));
 sky130_fd_sc_hd__xnor2_1 _14247_ (.A(_06915_),
    .B(_06917_),
    .Y(_06936_));
 sky130_fd_sc_hd__xor2_1 _14248_ (.A(_06935_),
    .B(_06936_),
    .X(_06937_));
 sky130_fd_sc_hd__nand2_1 _14249_ (.A(_06799_),
    .B(_06937_),
    .Y(_06938_));
 sky130_fd_sc_hd__o21a_1 _14250_ (.A1(_06935_),
    .A2(_06936_),
    .B1(_06938_),
    .X(_06939_));
 sky130_fd_sc_hd__or2_1 _14251_ (.A(_06933_),
    .B(_06939_),
    .X(_06940_));
 sky130_fd_sc_hd__or2_1 _14252_ (.A(_06921_),
    .B(_06929_),
    .X(_06941_));
 sky130_fd_sc_hd__nand2_1 _14253_ (.A(_06930_),
    .B(_06941_),
    .Y(_06942_));
 sky130_fd_sc_hd__nor2_1 _14254_ (.A(_06940_),
    .B(_06942_),
    .Y(_06943_));
 sky130_fd_sc_hd__nand2_1 _14255_ (.A(_06933_),
    .B(_06939_),
    .Y(_06944_));
 sky130_fd_sc_hd__or2_1 _14256_ (.A(_06799_),
    .B(_06937_),
    .X(_06945_));
 sky130_fd_sc_hd__nand2_1 _14257_ (.A(_06914_),
    .B(_06934_),
    .Y(_06946_));
 sky130_fd_sc_hd__inv_2 _14258_ (.A(_06934_),
    .Y(_06947_));
 sky130_fd_sc_hd__o211a_1 _14259_ (.A1(_06844_),
    .A2(_06914_),
    .B1(_06920_),
    .C1(_06947_),
    .X(_06948_));
 sky130_fd_sc_hd__a31o_1 _14260_ (.A1(_06844_),
    .A2(_06935_),
    .A3(_06946_),
    .B1(_06948_),
    .X(_06949_));
 sky130_fd_sc_hd__and4_1 _14261_ (.A(_06938_),
    .B(_06940_),
    .C(_06945_),
    .D(_06949_),
    .X(_06950_));
 sky130_fd_sc_hd__nand2_1 _14262_ (.A(_06940_),
    .B(_06942_),
    .Y(_06951_));
 sky130_fd_sc_hd__and4_1 _14263_ (.A(_06931_),
    .B(_06944_),
    .C(_06950_),
    .D(_06951_),
    .X(_06952_));
 sky130_fd_sc_hd__a21oi_1 _14264_ (.A1(_06927_),
    .A2(_06930_),
    .B1(_06908_),
    .Y(_06953_));
 sky130_fd_sc_hd__a211o_1 _14265_ (.A1(_06931_),
    .A2(_06943_),
    .B1(_06952_),
    .C1(_06953_),
    .X(_06954_));
 sky130_fd_sc_hd__nor2_1 _14266_ (.A(_06885_),
    .B(_06905_),
    .Y(_06955_));
 sky130_fd_sc_hd__a211o_1 _14267_ (.A1(_06906_),
    .A2(_06954_),
    .B1(_06955_),
    .C1(_06903_),
    .X(_06956_));
 sky130_fd_sc_hd__nor2_1 _14268_ (.A(_06875_),
    .B(_06874_),
    .Y(_06957_));
 sky130_fd_sc_hd__xnor2_1 _14269_ (.A(_06851_),
    .B(_06957_),
    .Y(_06958_));
 sky130_fd_sc_hd__and4_2 _14270_ (.A(_06879_),
    .B(_06880_),
    .C(_06956_),
    .D(_06958_),
    .X(_06959_));
 sky130_fd_sc_hd__a21oi_1 _14271_ (.A1(_06877_),
    .A2(_06879_),
    .B1(_06840_),
    .Y(_06960_));
 sky130_fd_sc_hd__xnor2_2 _14272_ (.A(_06795_),
    .B(_06960_),
    .Y(_06961_));
 sky130_fd_sc_hd__a32o_1 _14273_ (.A1(_06795_),
    .A2(_06877_),
    .A3(_06879_),
    .B1(_06959_),
    .B2(_06961_),
    .X(_06962_));
 sky130_fd_sc_hd__nor2_1 _14274_ (.A(_06782_),
    .B(_06841_),
    .Y(_06963_));
 sky130_fd_sc_hd__xnor2_1 _14275_ (.A(_06788_),
    .B(_06963_),
    .Y(_06964_));
 sky130_fd_sc_hd__and3_1 _14276_ (.A(_06790_),
    .B(_06782_),
    .C(_06788_),
    .X(_06965_));
 sky130_fd_sc_hd__a221o_1 _14277_ (.A1(_06788_),
    .A2(_06841_),
    .B1(_06962_),
    .B2(_06964_),
    .C1(_06965_),
    .X(_06966_));
 sky130_fd_sc_hd__xnor2_1 _14278_ (.A(_06686_),
    .B(_06688_),
    .Y(_06967_));
 sky130_fd_sc_hd__and2_1 _14279_ (.A(_06688_),
    .B(_06791_),
    .X(_06968_));
 sky130_fd_sc_hd__o21ba_1 _14280_ (.A1(_06791_),
    .A2(_06967_),
    .B1_N(_06968_),
    .X(_06969_));
 sky130_fd_sc_hd__a31o_1 _14281_ (.A1(_06794_),
    .A2(_06966_),
    .A3(_06969_),
    .B1(_06968_),
    .X(_06970_));
 sky130_fd_sc_hd__or2b_1 _14282_ (.A(_06631_),
    .B_N(_06689_),
    .X(_06971_));
 sky130_fd_sc_hd__a21oi_1 _14283_ (.A1(_06629_),
    .A2(_06971_),
    .B1(_06573_),
    .Y(_06972_));
 sky130_fd_sc_hd__a31o_1 _14284_ (.A1(_06630_),
    .A2(_06690_),
    .A3(_06970_),
    .B1(_06972_),
    .X(_06973_));
 sky130_fd_sc_hd__a211o_1 _14285_ (.A1(_06571_),
    .A2(_06973_),
    .B1(_06567_),
    .C1(_06569_),
    .X(_06974_));
 sky130_fd_sc_hd__nand2_1 _14286_ (.A(_06455_),
    .B(_06974_),
    .Y(_06975_));
 sky130_fd_sc_hd__or3b_1 _14287_ (.A(_06372_),
    .B(_06399_),
    .C_N(_06401_),
    .X(_06976_));
 sky130_fd_sc_hd__o21ai_1 _14288_ (.A1(_06453_),
    .A2(_06402_),
    .B1(_06976_),
    .Y(_06977_));
 sky130_fd_sc_hd__nand2_1 _14289_ (.A(_06370_),
    .B(_06977_),
    .Y(_06978_));
 sky130_fd_sc_hd__o31a_2 _14290_ (.A1(_06371_),
    .A2(_06402_),
    .A3(_06975_),
    .B1(_06978_),
    .X(_06979_));
 sky130_fd_sc_hd__xor2_2 _14291_ (.A(_06368_),
    .B(_06979_),
    .X(_06980_));
 sky130_fd_sc_hd__buf_2 _14292_ (.A(_05593_),
    .X(_06981_));
 sky130_fd_sc_hd__a21boi_1 _14293_ (.A1(_06455_),
    .A2(_06974_),
    .B1_N(_06453_),
    .Y(_06982_));
 sky130_fd_sc_hd__o211ai_1 _14294_ (.A1(_06402_),
    .A2(_06982_),
    .B1(_06976_),
    .C1(_06371_),
    .Y(_06983_));
 sky130_fd_sc_hd__and3_1 _14295_ (.A(_06981_),
    .B(_06979_),
    .C(_06983_),
    .X(_06984_));
 sky130_fd_sc_hd__buf_2 _14296_ (.A(_05501_),
    .X(_06985_));
 sky130_fd_sc_hd__a211o_1 _14297_ (.A1(_05432_),
    .A2(_06980_),
    .B1(_06984_),
    .C1(_06985_),
    .X(_06986_));
 sky130_fd_sc_hd__buf_2 _14298_ (.A(_05586_),
    .X(_06987_));
 sky130_fd_sc_hd__or3_1 _14299_ (.A(_05432_),
    .B(_06368_),
    .C(_06979_),
    .X(_06988_));
 sky130_fd_sc_hd__or3b_1 _14300_ (.A(_05434_),
    .B(_06987_),
    .C_N(_06988_),
    .X(_06989_));
 sky130_fd_sc_hd__buf_2 _14301_ (.A(_05531_),
    .X(_06990_));
 sky130_fd_sc_hd__a21o_1 _14302_ (.A1(_06986_),
    .A2(_06989_),
    .B1(_06990_),
    .X(_06991_));
 sky130_fd_sc_hd__xor2_1 _14303_ (.A(_06402_),
    .B(_06982_),
    .X(_06992_));
 sky130_fd_sc_hd__xor2_1 _14304_ (.A(_06455_),
    .B(_06974_),
    .X(_06993_));
 sky130_fd_sc_hd__and2_1 _14305_ (.A(_06981_),
    .B(_06993_),
    .X(_06994_));
 sky130_fd_sc_hd__a21o_1 _14306_ (.A1(_05432_),
    .A2(_06992_),
    .B1(_06994_),
    .X(_06995_));
 sky130_fd_sc_hd__xor2_1 _14307_ (.A(_06571_),
    .B(_06973_),
    .X(_06996_));
 sky130_fd_sc_hd__and2_1 _14308_ (.A(_05431_),
    .B(_06996_),
    .X(_06997_));
 sky130_fd_sc_hd__or2_1 _14309_ (.A(_06573_),
    .B(_06629_),
    .X(_06998_));
 sky130_fd_sc_hd__and2_1 _14310_ (.A(_06630_),
    .B(_06998_),
    .X(_06999_));
 sky130_fd_sc_hd__a21boi_1 _14311_ (.A1(_06690_),
    .A2(_06970_),
    .B1_N(_06971_),
    .Y(_07000_));
 sky130_fd_sc_hd__xnor2_1 _14312_ (.A(_06999_),
    .B(_07000_),
    .Y(_07001_));
 sky130_fd_sc_hd__and2_1 _14313_ (.A(_05593_),
    .B(_07001_),
    .X(_07002_));
 sky130_fd_sc_hd__or2_1 _14314_ (.A(_06997_),
    .B(_07002_),
    .X(_07003_));
 sky130_fd_sc_hd__or2_1 _14315_ (.A(_06985_),
    .B(_07003_),
    .X(_07004_));
 sky130_fd_sc_hd__o21ai_1 _14316_ (.A1(_06987_),
    .A2(_06995_),
    .B1(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__nand2_1 _14317_ (.A(_06990_),
    .B(_07005_),
    .Y(_07006_));
 sky130_fd_sc_hd__clkbuf_2 _14318_ (.A(_05569_),
    .X(_07007_));
 sky130_fd_sc_hd__and2_1 _14319_ (.A(_06962_),
    .B(_06964_),
    .X(_07008_));
 sky130_fd_sc_hd__nor2_1 _14320_ (.A(_06962_),
    .B(_06964_),
    .Y(_07009_));
 sky130_fd_sc_hd__or2_1 _14321_ (.A(_07008_),
    .B(_07009_),
    .X(_07010_));
 sky130_fd_sc_hd__nor2_1 _14322_ (.A(_05431_),
    .B(_07010_),
    .Y(_07011_));
 sky130_fd_sc_hd__a21oi_1 _14323_ (.A1(_06788_),
    .A2(_06841_),
    .B1(_07008_),
    .Y(_07012_));
 sky130_fd_sc_hd__o21ba_1 _14324_ (.A1(_06789_),
    .A2(_06793_),
    .B1_N(_06965_),
    .X(_07013_));
 sky130_fd_sc_hd__xnor2_1 _14325_ (.A(_07012_),
    .B(_07013_),
    .Y(_07014_));
 sky130_fd_sc_hd__and2_1 _14326_ (.A(_05431_),
    .B(_07014_),
    .X(_07015_));
 sky130_fd_sc_hd__or2_1 _14327_ (.A(_07011_),
    .B(_07015_),
    .X(_07016_));
 sky130_fd_sc_hd__xor2_1 _14328_ (.A(_06690_),
    .B(_06970_),
    .X(_07017_));
 sky130_fd_sc_hd__and2_1 _14329_ (.A(_05431_),
    .B(_07017_),
    .X(_07018_));
 sky130_fd_sc_hd__nand2_1 _14330_ (.A(_06794_),
    .B(_06966_),
    .Y(_07019_));
 sky130_fd_sc_hd__xnor2_1 _14331_ (.A(_07019_),
    .B(_06969_),
    .Y(_07020_));
 sky130_fd_sc_hd__nand2_1 _14332_ (.A(_06981_),
    .B(_07020_),
    .Y(_07021_));
 sky130_fd_sc_hd__or2b_1 _14333_ (.A(_07018_),
    .B_N(_07021_),
    .X(_07022_));
 sky130_fd_sc_hd__mux2_1 _14334_ (.A0(_07016_),
    .A1(_07022_),
    .S(_06985_),
    .X(_07023_));
 sky130_fd_sc_hd__xnor2_4 _14335_ (.A(_06959_),
    .B(_06961_),
    .Y(_07024_));
 sky130_fd_sc_hd__nor2_1 _14336_ (.A(_05515_),
    .B(_07024_),
    .Y(_07025_));
 sky130_fd_sc_hd__mux2_1 _14337_ (.A0(_07023_),
    .A1(_07025_),
    .S(_05531_),
    .X(_07026_));
 sky130_fd_sc_hd__and2_1 _14338_ (.A(_07007_),
    .B(_07026_),
    .X(_07027_));
 sky130_fd_sc_hd__a31oi_4 _14339_ (.A1(_05408_),
    .A2(_06991_),
    .A3(_07006_),
    .B1(_07027_),
    .Y(_07028_));
 sky130_fd_sc_hd__buf_2 _14340_ (.A(_05458_),
    .X(_07029_));
 sky130_fd_sc_hd__nor3_2 _14341_ (.A(_06981_),
    .B(_06368_),
    .C(_06979_),
    .Y(_07030_));
 sky130_fd_sc_hd__a21o_1 _14342_ (.A1(_06981_),
    .A2(_06980_),
    .B1(_07030_),
    .X(_07031_));
 sky130_fd_sc_hd__and2_1 _14343_ (.A(_06981_),
    .B(_06992_),
    .X(_07032_));
 sky130_fd_sc_hd__and3_1 _14344_ (.A(_05432_),
    .B(_06979_),
    .C(_06983_),
    .X(_07033_));
 sky130_fd_sc_hd__and2_1 _14345_ (.A(_06981_),
    .B(_06996_),
    .X(_07034_));
 sky130_fd_sc_hd__a21o_1 _14346_ (.A1(_05432_),
    .A2(_06993_),
    .B1(_07034_),
    .X(_07035_));
 sky130_fd_sc_hd__or2_1 _14347_ (.A(_06985_),
    .B(_07035_),
    .X(_07036_));
 sky130_fd_sc_hd__o311a_1 _14348_ (.A1(_06987_),
    .A2(_07032_),
    .A3(_07033_),
    .B1(_07036_),
    .C1(_06990_),
    .X(_07037_));
 sky130_fd_sc_hd__a31o_1 _14349_ (.A1(_07029_),
    .A2(_06987_),
    .A3(_07031_),
    .B1(_07037_),
    .X(_07038_));
 sky130_fd_sc_hd__and2_1 _14350_ (.A(_05593_),
    .B(_07014_),
    .X(_07039_));
 sky130_fd_sc_hd__nand2_1 _14351_ (.A(_05431_),
    .B(_07020_),
    .Y(_07040_));
 sky130_fd_sc_hd__or2b_1 _14352_ (.A(_07039_),
    .B_N(_07040_),
    .X(_07041_));
 sky130_fd_sc_hd__and2_1 _14353_ (.A(_06981_),
    .B(_07017_),
    .X(_07042_));
 sky130_fd_sc_hd__and2_1 _14354_ (.A(_05432_),
    .B(_07001_),
    .X(_07043_));
 sky130_fd_sc_hd__or3_1 _14355_ (.A(_05586_),
    .B(_07042_),
    .C(_07043_),
    .X(_07044_));
 sky130_fd_sc_hd__o21a_1 _14356_ (.A1(_06985_),
    .A2(_07041_),
    .B1(_07044_),
    .X(_07045_));
 sky130_fd_sc_hd__nor2_1 _14357_ (.A(_05431_),
    .B(_07024_),
    .Y(_07046_));
 sky130_fd_sc_hd__nor2_1 _14358_ (.A(_05593_),
    .B(_07010_),
    .Y(_07047_));
 sky130_fd_sc_hd__nor2_1 _14359_ (.A(_07046_),
    .B(_07047_),
    .Y(_07048_));
 sky130_fd_sc_hd__nor2_1 _14360_ (.A(_06987_),
    .B(_07048_),
    .Y(_07049_));
 sky130_fd_sc_hd__mux2_1 _14361_ (.A0(_07045_),
    .A1(_07049_),
    .S(_05531_),
    .X(_07050_));
 sky130_fd_sc_hd__or2_1 _14362_ (.A(_05408_),
    .B(_07050_),
    .X(_07051_));
 sky130_fd_sc_hd__o21ai_1 _14363_ (.A1(_07007_),
    .A2(_07038_),
    .B1(_07051_),
    .Y(_07052_));
 sky130_fd_sc_hd__or2_1 _14364_ (.A(_06985_),
    .B(_06995_),
    .X(_07053_));
 sky130_fd_sc_hd__a211o_1 _14365_ (.A1(_05432_),
    .A2(_06980_),
    .B1(_06984_),
    .C1(_06987_),
    .X(_07054_));
 sky130_fd_sc_hd__mux2_1 _14366_ (.A0(_07003_),
    .A1(_07022_),
    .S(_05586_),
    .X(_07055_));
 sky130_fd_sc_hd__and2_1 _14367_ (.A(_05531_),
    .B(_07055_),
    .X(_07056_));
 sky130_fd_sc_hd__a31o_1 _14368_ (.A1(_07029_),
    .A2(_07053_),
    .A3(_07054_),
    .B1(_07056_),
    .X(_07057_));
 sky130_fd_sc_hd__or2_1 _14369_ (.A(_05593_),
    .B(_07024_),
    .X(_07058_));
 sky130_fd_sc_hd__inv_2 _14370_ (.A(_07058_),
    .Y(_07059_));
 sky130_fd_sc_hd__mux2_1 _14371_ (.A0(_07016_),
    .A1(_07059_),
    .S(_05586_),
    .X(_07060_));
 sky130_fd_sc_hd__nand2_1 _14372_ (.A(_07029_),
    .B(_07060_),
    .Y(_07061_));
 sky130_fd_sc_hd__nor2_1 _14373_ (.A(_05408_),
    .B(_07061_),
    .Y(_07062_));
 sky130_fd_sc_hd__a21oi_1 _14374_ (.A1(_05408_),
    .A2(_07057_),
    .B1(_07062_),
    .Y(_07063_));
 sky130_fd_sc_hd__a211o_1 _14375_ (.A1(_06981_),
    .A2(_06980_),
    .B1(_07030_),
    .C1(_06987_),
    .X(_07064_));
 sky130_fd_sc_hd__or3_1 _14376_ (.A(_06985_),
    .B(_07032_),
    .C(_07033_),
    .X(_07065_));
 sky130_fd_sc_hd__or3_1 _14377_ (.A(_05501_),
    .B(_07042_),
    .C(_07043_),
    .X(_07066_));
 sky130_fd_sc_hd__o21ai_1 _14378_ (.A1(_05586_),
    .A2(_07035_),
    .B1(_07066_),
    .Y(_07067_));
 sky130_fd_sc_hd__nor2_1 _14379_ (.A(_07029_),
    .B(_07067_),
    .Y(_07068_));
 sky130_fd_sc_hd__a31o_1 _14380_ (.A1(_07029_),
    .A2(_07064_),
    .A3(_07065_),
    .B1(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__clkinv_2 _14381_ (.A(_07048_),
    .Y(_07070_));
 sky130_fd_sc_hd__mux2_1 _14382_ (.A0(_07041_),
    .A1(_07070_),
    .S(_05586_),
    .X(_07071_));
 sky130_fd_sc_hd__nand2_1 _14383_ (.A(_07029_),
    .B(_07071_),
    .Y(_07072_));
 sky130_fd_sc_hd__nor2_1 _14384_ (.A(_05408_),
    .B(_07072_),
    .Y(_07073_));
 sky130_fd_sc_hd__a21oi_1 _14385_ (.A1(_05408_),
    .A2(_07069_),
    .B1(_07073_),
    .Y(_07074_));
 sky130_fd_sc_hd__or2_2 _14386_ (.A(_05440_),
    .B(_05405_),
    .X(_07075_));
 sky130_fd_sc_hd__a41o_1 _14387_ (.A1(_07028_),
    .A2(_07052_),
    .A3(_07063_),
    .A4(_07074_),
    .B1(_07075_),
    .X(_07076_));
 sky130_fd_sc_hd__o311a_1 _14388_ (.A1(_06987_),
    .A2(_07032_),
    .A3(_07033_),
    .B1(_07036_),
    .C1(_07029_),
    .X(_07077_));
 sky130_fd_sc_hd__a21oi_1 _14389_ (.A1(_06990_),
    .A2(_07045_),
    .B1(_07077_),
    .Y(_07078_));
 sky130_fd_sc_hd__and2_1 _14390_ (.A(_07029_),
    .B(_05404_),
    .X(_07079_));
 sky130_fd_sc_hd__a2bb2o_1 _14391_ (.A1_N(_07007_),
    .A2_N(_07078_),
    .B1(_07079_),
    .B2(_07049_),
    .X(_07080_));
 sky130_fd_sc_hd__clkinv_2 _14392_ (.A(_07023_),
    .Y(_07081_));
 sky130_fd_sc_hd__mux2_1 _14393_ (.A0(_07005_),
    .A1(_07081_),
    .S(_06990_),
    .X(_07082_));
 sky130_fd_sc_hd__a2bb2o_1 _14394_ (.A1_N(_07007_),
    .A2_N(_07082_),
    .B1(_07079_),
    .B2(_07025_),
    .X(_07083_));
 sky130_fd_sc_hd__inv_2 _14395_ (.A(_07071_),
    .Y(_07084_));
 sky130_fd_sc_hd__mux2_1 _14396_ (.A0(_07067_),
    .A1(_07084_),
    .S(_05531_),
    .X(_07085_));
 sky130_fd_sc_hd__nor2_1 _14397_ (.A(_05569_),
    .B(_07085_),
    .Y(_07086_));
 sky130_fd_sc_hd__or2_1 _14398_ (.A(_07029_),
    .B(_07060_),
    .X(_07087_));
 sky130_fd_sc_hd__o21ai_1 _14399_ (.A1(_05531_),
    .A2(_07055_),
    .B1(_07087_),
    .Y(_07088_));
 sky130_fd_sc_hd__or2_1 _14400_ (.A(_05569_),
    .B(_07088_),
    .X(_07089_));
 sky130_fd_sc_hd__or3b_1 _14401_ (.A(_07075_),
    .B(_07086_),
    .C_N(_07089_),
    .X(_07090_));
 sky130_fd_sc_hd__a211oi_1 _14402_ (.A1(_05401_),
    .A2(_06988_),
    .B1(_06985_),
    .C1(_05531_),
    .Y(_07091_));
 sky130_fd_sc_hd__a31o_1 _14403_ (.A1(_06990_),
    .A2(_07053_),
    .A3(_07054_),
    .B1(_07091_),
    .X(_07092_));
 sky130_fd_sc_hd__and3_1 _14404_ (.A(_06990_),
    .B(_06986_),
    .C(_06989_),
    .X(_07093_));
 sky130_fd_sc_hd__and3_1 _14405_ (.A(_06990_),
    .B(_07064_),
    .C(_07065_),
    .X(_07094_));
 sky130_fd_sc_hd__a31o_1 _14406_ (.A1(_06990_),
    .A2(_06987_),
    .A3(_07031_),
    .B1(_05568_),
    .X(_07095_));
 sky130_fd_sc_hd__nand2_1 _14407_ (.A(_07075_),
    .B(_05408_),
    .Y(_07096_));
 sky130_fd_sc_hd__o41a_1 _14408_ (.A1(_07092_),
    .A2(_07093_),
    .A3(_07094_),
    .A4(_07095_),
    .B1(_07096_),
    .X(_07097_));
 sky130_fd_sc_hd__o31ai_4 _14409_ (.A1(_07080_),
    .A2(_07083_),
    .A3(_07090_),
    .B1(_07097_),
    .Y(_07098_));
 sky130_fd_sc_hd__a21o_2 _14410_ (.A1(_07076_),
    .A2(_07098_),
    .B1(_05538_),
    .X(_07099_));
 sky130_fd_sc_hd__clkbuf_4 _14411_ (.A(_07099_),
    .X(_07100_));
 sky130_fd_sc_hd__clkbuf_4 _14412_ (.A(_07100_),
    .X(_07101_));
 sky130_fd_sc_hd__buf_4 _14413_ (.A(_07101_),
    .X(_07102_));
 sky130_fd_sc_hd__or2_1 _14414_ (.A(_06997_),
    .B(_06994_),
    .X(_07103_));
 sky130_fd_sc_hd__a21o_1 _14415_ (.A1(_05432_),
    .A2(_06992_),
    .B1(_06984_),
    .X(_07104_));
 sky130_fd_sc_hd__buf_2 _14416_ (.A(_05497_),
    .X(_07105_));
 sky130_fd_sc_hd__mux2_1 _14417_ (.A0(_07103_),
    .A1(_07104_),
    .S(_07105_),
    .X(_07106_));
 sky130_fd_sc_hd__buf_2 _14418_ (.A(_05499_),
    .X(_07107_));
 sky130_fd_sc_hd__a21bo_1 _14419_ (.A1(_05432_),
    .A2(_06980_),
    .B1_N(_06988_),
    .X(_07108_));
 sky130_fd_sc_hd__and3_1 _14420_ (.A(_05517_),
    .B(_07107_),
    .C(_07108_),
    .X(_07109_));
 sky130_fd_sc_hd__a21oi_1 _14421_ (.A1(_05527_),
    .A2(_07106_),
    .B1(_07109_),
    .Y(_07110_));
 sky130_fd_sc_hd__or2b_1 _14422_ (.A(_07015_),
    .B_N(_07021_),
    .X(_07111_));
 sky130_fd_sc_hd__or2_1 _14423_ (.A(_07002_),
    .B(_07018_),
    .X(_07112_));
 sky130_fd_sc_hd__mux2_1 _14424_ (.A0(_07111_),
    .A1(_07112_),
    .S(_07105_),
    .X(_07113_));
 sky130_fd_sc_hd__or2_1 _14425_ (.A(_07011_),
    .B(_07059_),
    .X(_07114_));
 sky130_fd_sc_hd__nor2_1 _14426_ (.A(_05517_),
    .B(_05499_),
    .Y(_07115_));
 sky130_fd_sc_hd__a221oi_1 _14427_ (.A1(_07107_),
    .A2(_07113_),
    .B1(_07114_),
    .B2(_07115_),
    .C1(_05577_),
    .Y(_07116_));
 sky130_fd_sc_hd__a211o_1 _14428_ (.A1(_05577_),
    .A2(_07110_),
    .B1(_07116_),
    .C1(_05602_),
    .X(_07117_));
 sky130_fd_sc_hd__nand2_1 _14429_ (.A(_07102_),
    .B(_07117_),
    .Y(_07118_));
 sky130_fd_sc_hd__mux2_1 _14430_ (.A0(\rbzero.wall_tracer.stepDistY[-12] ),
    .A1(_07118_),
    .S(_00004_),
    .X(_07119_));
 sky130_fd_sc_hd__clkbuf_1 _14431_ (.A(_07119_),
    .X(_00406_));
 sky130_fd_sc_hd__a21oi_1 _14432_ (.A1(_05432_),
    .A2(_06993_),
    .B1(_07032_),
    .Y(_07120_));
 sky130_fd_sc_hd__a21o_1 _14433_ (.A1(_06981_),
    .A2(_06980_),
    .B1(_07033_),
    .X(_07121_));
 sky130_fd_sc_hd__nand2_1 _14434_ (.A(_07105_),
    .B(_07121_),
    .Y(_07122_));
 sky130_fd_sc_hd__o21a_1 _14435_ (.A1(_07105_),
    .A2(_07120_),
    .B1(_07122_),
    .X(_07123_));
 sky130_fd_sc_hd__o32a_1 _14436_ (.A1(_05459_),
    .A2(_06368_),
    .A3(_06979_),
    .B1(_07123_),
    .B2(_07107_),
    .X(_07124_));
 sky130_fd_sc_hd__and2b_1 _14437_ (.A_N(_07042_),
    .B(_07040_),
    .X(_07125_));
 sky130_fd_sc_hd__or2_1 _14438_ (.A(_07105_),
    .B(_07125_),
    .X(_07126_));
 sky130_fd_sc_hd__nor2_1 _14439_ (.A(_07043_),
    .B(_07034_),
    .Y(_07127_));
 sky130_fd_sc_hd__or2_1 _14440_ (.A(_05517_),
    .B(_07127_),
    .X(_07128_));
 sky130_fd_sc_hd__a21oi_1 _14441_ (.A1(_07126_),
    .A2(_07128_),
    .B1(_05527_),
    .Y(_07129_));
 sky130_fd_sc_hd__nor2_1 _14442_ (.A(_07105_),
    .B(_05499_),
    .Y(_07130_));
 sky130_fd_sc_hd__or2_1 _14443_ (.A(_07039_),
    .B(_07047_),
    .X(_07131_));
 sky130_fd_sc_hd__a22o_1 _14444_ (.A1(_07130_),
    .A2(_07046_),
    .B1(_07131_),
    .B2(_07115_),
    .X(_07132_));
 sky130_fd_sc_hd__clkbuf_4 _14445_ (.A(_05538_),
    .X(_07133_));
 sky130_fd_sc_hd__o31a_1 _14446_ (.A1(_05577_),
    .A2(_07129_),
    .A3(_07132_),
    .B1(_07133_),
    .X(_07134_));
 sky130_fd_sc_hd__a21bo_1 _14447_ (.A1(_05577_),
    .A2(_07124_),
    .B1_N(_07134_),
    .X(_07135_));
 sky130_fd_sc_hd__nand2_1 _14448_ (.A(_07102_),
    .B(_07135_),
    .Y(_07136_));
 sky130_fd_sc_hd__mux2_1 _14449_ (.A0(\rbzero.wall_tracer.stepDistY[-11] ),
    .A1(_07136_),
    .S(_00004_),
    .X(_07137_));
 sky130_fd_sc_hd__clkbuf_1 _14450_ (.A(_07137_),
    .X(_00407_));
 sky130_fd_sc_hd__or2_1 _14451_ (.A(_05497_),
    .B(_07104_),
    .X(_07138_));
 sky130_fd_sc_hd__o21ai_1 _14452_ (.A1(_05517_),
    .A2(_07108_),
    .B1(_07138_),
    .Y(_07139_));
 sky130_fd_sc_hd__o21a_1 _14453_ (.A1(_07107_),
    .A2(_07139_),
    .B1(_05401_),
    .X(_07140_));
 sky130_fd_sc_hd__nand2_1 _14454_ (.A(_05517_),
    .B(_07112_),
    .Y(_07141_));
 sky130_fd_sc_hd__nand2_1 _14455_ (.A(_07105_),
    .B(_07103_),
    .Y(_07142_));
 sky130_fd_sc_hd__a21oi_1 _14456_ (.A1(_07141_),
    .A2(_07142_),
    .B1(_05527_),
    .Y(_07143_));
 sky130_fd_sc_hd__a22o_1 _14457_ (.A1(_07115_),
    .A2(_07111_),
    .B1(_07114_),
    .B2(_07130_),
    .X(_07144_));
 sky130_fd_sc_hd__o31ai_1 _14458_ (.A1(_05577_),
    .A2(_07143_),
    .A3(_07144_),
    .B1(_07133_),
    .Y(_07145_));
 sky130_fd_sc_hd__a21o_1 _14459_ (.A1(_05577_),
    .A2(_07140_),
    .B1(_07145_),
    .X(_07146_));
 sky130_fd_sc_hd__nand2_1 _14460_ (.A(_07102_),
    .B(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__mux2_1 _14461_ (.A0(\rbzero.wall_tracer.stepDistY[-10] ),
    .A1(_07147_),
    .S(_00004_),
    .X(_07148_));
 sky130_fd_sc_hd__clkbuf_1 _14462_ (.A(_07148_),
    .X(_00408_));
 sky130_fd_sc_hd__a22oi_1 _14463_ (.A1(_06987_),
    .A2(_07030_),
    .B1(_07121_),
    .B2(_05517_),
    .Y(_07149_));
 sky130_fd_sc_hd__or2_1 _14464_ (.A(_07107_),
    .B(_07149_),
    .X(_07150_));
 sky130_fd_sc_hd__mux2_1 _14465_ (.A0(_07127_),
    .A1(_07120_),
    .S(_07105_),
    .X(_07151_));
 sky130_fd_sc_hd__nor2_1 _14466_ (.A(_07105_),
    .B(_07131_),
    .Y(_07152_));
 sky130_fd_sc_hd__a211o_1 _14467_ (.A1(_07105_),
    .A2(_07125_),
    .B1(_07152_),
    .C1(_07107_),
    .X(_07153_));
 sky130_fd_sc_hd__o211a_1 _14468_ (.A1(_05527_),
    .A2(_07151_),
    .B1(_07153_),
    .C1(_05535_),
    .X(_07154_));
 sky130_fd_sc_hd__a211oi_1 _14469_ (.A1(_05577_),
    .A2(_07150_),
    .B1(_07154_),
    .C1(_05602_),
    .Y(_07155_));
 sky130_fd_sc_hd__a21oi_2 _14470_ (.A1(_05470_),
    .A2(_07049_),
    .B1(_07155_),
    .Y(_07156_));
 sky130_fd_sc_hd__nand2_1 _14471_ (.A(_07102_),
    .B(_07156_),
    .Y(_07157_));
 sky130_fd_sc_hd__mux2_1 _14472_ (.A0(\rbzero.wall_tracer.stepDistY[-9] ),
    .A1(_07157_),
    .S(_00004_),
    .X(_07158_));
 sky130_fd_sc_hd__clkbuf_1 _14473_ (.A(_07158_),
    .X(_00409_));
 sky130_fd_sc_hd__nand2_1 _14474_ (.A(_05602_),
    .B(_05408_),
    .Y(_07159_));
 sky130_fd_sc_hd__a21o_1 _14475_ (.A1(_05527_),
    .A2(_07113_),
    .B1(_05577_),
    .X(_07160_));
 sky130_fd_sc_hd__a21oi_1 _14476_ (.A1(_07107_),
    .A2(_07106_),
    .B1(_07160_),
    .Y(_07161_));
 sky130_fd_sc_hd__nand2_2 _14477_ (.A(_07130_),
    .B(_07108_),
    .Y(_07162_));
 sky130_fd_sc_hd__a21o_1 _14478_ (.A1(_05447_),
    .A2(_07162_),
    .B1(_05602_),
    .X(_07163_));
 sky130_fd_sc_hd__o22a_2 _14479_ (.A1(_07159_),
    .A2(_07061_),
    .B1(_07161_),
    .B2(_07163_),
    .X(_07164_));
 sky130_fd_sc_hd__nand2_2 _14480_ (.A(_07102_),
    .B(_07164_),
    .Y(_07165_));
 sky130_fd_sc_hd__mux2_1 _14481_ (.A0(\rbzero.wall_tracer.stepDistY[-8] ),
    .A1(_07165_),
    .S(_00004_),
    .X(_07166_));
 sky130_fd_sc_hd__clkbuf_1 _14482_ (.A(_07166_),
    .X(_00410_));
 sky130_fd_sc_hd__a21o_1 _14483_ (.A1(_07126_),
    .A2(_07128_),
    .B1(_07107_),
    .X(_07167_));
 sky130_fd_sc_hd__o211a_1 _14484_ (.A1(_05527_),
    .A2(_07123_),
    .B1(_07167_),
    .C1(_05535_),
    .X(_07168_));
 sky130_fd_sc_hd__nand2_1 _14485_ (.A(_07130_),
    .B(_07030_),
    .Y(_07169_));
 sky130_fd_sc_hd__a21o_1 _14486_ (.A1(_05447_),
    .A2(_07169_),
    .B1(_05602_),
    .X(_07170_));
 sky130_fd_sc_hd__o22a_2 _14487_ (.A1(_07159_),
    .A2(_07072_),
    .B1(_07168_),
    .B2(_07170_),
    .X(_07171_));
 sky130_fd_sc_hd__nand2_2 _14488_ (.A(_07102_),
    .B(_07171_),
    .Y(_07172_));
 sky130_fd_sc_hd__mux2_1 _14489_ (.A0(\rbzero.wall_tracer.stepDistY[-7] ),
    .A1(_07172_),
    .S(_00004_),
    .X(_07173_));
 sky130_fd_sc_hd__clkbuf_1 _14490_ (.A(_07173_),
    .X(_00411_));
 sky130_fd_sc_hd__nor2_1 _14491_ (.A(_07133_),
    .B(_07007_),
    .Y(_07174_));
 sky130_fd_sc_hd__and3_1 _14492_ (.A(_05527_),
    .B(_07141_),
    .C(_07142_),
    .X(_07175_));
 sky130_fd_sc_hd__or2_1 _14493_ (.A(_05602_),
    .B(_05577_),
    .X(_07176_));
 sky130_fd_sc_hd__buf_2 _14494_ (.A(_07176_),
    .X(_07177_));
 sky130_fd_sc_hd__a21o_1 _14495_ (.A1(_07107_),
    .A2(_07139_),
    .B1(_07177_),
    .X(_07178_));
 sky130_fd_sc_hd__o2bb2a_2 _14496_ (.A1_N(_07174_),
    .A2_N(_07026_),
    .B1(_07175_),
    .B2(_07178_),
    .X(_07179_));
 sky130_fd_sc_hd__nand2_2 _14497_ (.A(_07102_),
    .B(_07179_),
    .Y(_07180_));
 sky130_fd_sc_hd__mux2_1 _14498_ (.A0(\rbzero.wall_tracer.stepDistY[-6] ),
    .A1(_07180_),
    .S(_00004_),
    .X(_07181_));
 sky130_fd_sc_hd__clkbuf_1 _14499_ (.A(_07181_),
    .X(_00412_));
 sky130_fd_sc_hd__a21o_1 _14500_ (.A1(_05527_),
    .A2(_07151_),
    .B1(_07177_),
    .X(_07182_));
 sky130_fd_sc_hd__a21oi_1 _14501_ (.A1(_07107_),
    .A2(_07149_),
    .B1(_07182_),
    .Y(_07183_));
 sky130_fd_sc_hd__a21oi_4 _14502_ (.A1(_07174_),
    .A2(_07050_),
    .B1(_07183_),
    .Y(_07184_));
 sky130_fd_sc_hd__nand2_2 _14503_ (.A(_07102_),
    .B(_07184_),
    .Y(_07185_));
 sky130_fd_sc_hd__mux2_1 _14504_ (.A0(\rbzero.wall_tracer.stepDistY[-5] ),
    .A1(_07185_),
    .S(_00004_),
    .X(_07186_));
 sky130_fd_sc_hd__clkbuf_1 _14505_ (.A(_07186_),
    .X(_00413_));
 sky130_fd_sc_hd__or2_1 _14506_ (.A(_07177_),
    .B(_07110_),
    .X(_07187_));
 sky130_fd_sc_hd__or2_1 _14507_ (.A(_07133_),
    .B(_07089_),
    .X(_07188_));
 sky130_fd_sc_hd__nand3_4 _14508_ (.A(_07101_),
    .B(_07187_),
    .C(_07188_),
    .Y(_07189_));
 sky130_fd_sc_hd__mux2_1 _14509_ (.A0(\rbzero.wall_tracer.stepDistY[-4] ),
    .A1(_07189_),
    .S(_00004_),
    .X(_07190_));
 sky130_fd_sc_hd__clkbuf_1 _14510_ (.A(_07190_),
    .X(_00414_));
 sky130_fd_sc_hd__o2bb2a_1 _14511_ (.A1_N(_05602_),
    .A2_N(_07086_),
    .B1(_07124_),
    .B2(_07177_),
    .X(_07191_));
 sky130_fd_sc_hd__nand2_1 _14512_ (.A(_07102_),
    .B(_07191_),
    .Y(_07192_));
 sky130_fd_sc_hd__clkbuf_4 _14513_ (.A(_04925_),
    .X(_07193_));
 sky130_fd_sc_hd__mux2_1 _14514_ (.A0(\rbzero.wall_tracer.stepDistY[-3] ),
    .A1(_07192_),
    .S(_07193_),
    .X(_07194_));
 sky130_fd_sc_hd__clkbuf_1 _14515_ (.A(_07194_),
    .X(_00415_));
 sky130_fd_sc_hd__o2bb2a_2 _14516_ (.A1_N(_05602_),
    .A2_N(_07083_),
    .B1(_07140_),
    .B2(_07177_),
    .X(_07195_));
 sky130_fd_sc_hd__nand2_1 _14517_ (.A(_07102_),
    .B(_07195_),
    .Y(_07196_));
 sky130_fd_sc_hd__mux2_1 _14518_ (.A0(\rbzero.wall_tracer.stepDistY[-2] ),
    .A1(_07196_),
    .S(_07193_),
    .X(_07197_));
 sky130_fd_sc_hd__clkbuf_1 _14519_ (.A(_07197_),
    .X(_00416_));
 sky130_fd_sc_hd__o2bb2a_1 _14520_ (.A1_N(_05602_),
    .A2_N(_07080_),
    .B1(_07150_),
    .B2(_07177_),
    .X(_07198_));
 sky130_fd_sc_hd__nand2_2 _14521_ (.A(_07101_),
    .B(_07198_),
    .Y(_07199_));
 sky130_fd_sc_hd__mux2_1 _14522_ (.A0(\rbzero.wall_tracer.stepDistY[-1] ),
    .A1(_07199_),
    .S(_07193_),
    .X(_07200_));
 sky130_fd_sc_hd__clkbuf_1 _14523_ (.A(_07200_),
    .X(_00417_));
 sky130_fd_sc_hd__or2_1 _14524_ (.A(_07133_),
    .B(_07063_),
    .X(_07201_));
 sky130_fd_sc_hd__o211ai_4 _14525_ (.A1(_07177_),
    .A2(_07162_),
    .B1(_07201_),
    .C1(_07099_),
    .Y(_07202_));
 sky130_fd_sc_hd__mux2_1 _14526_ (.A0(\rbzero.wall_tracer.stepDistY[0] ),
    .A1(_07202_),
    .S(_07193_),
    .X(_07203_));
 sky130_fd_sc_hd__clkbuf_1 _14527_ (.A(_07203_),
    .X(_00418_));
 sky130_fd_sc_hd__or2_1 _14528_ (.A(_07133_),
    .B(_07074_),
    .X(_07204_));
 sky130_fd_sc_hd__or2_1 _14529_ (.A(_07177_),
    .B(_07169_),
    .X(_07205_));
 sky130_fd_sc_hd__nand3_4 _14530_ (.A(_07099_),
    .B(_07204_),
    .C(_07205_),
    .Y(_07206_));
 sky130_fd_sc_hd__mux2_1 _14531_ (.A0(\rbzero.wall_tracer.stepDistY[1] ),
    .A1(_07206_),
    .S(_07193_),
    .X(_07207_));
 sky130_fd_sc_hd__clkbuf_1 _14532_ (.A(_07207_),
    .X(_00419_));
 sky130_fd_sc_hd__a31oi_4 _14533_ (.A1(_07028_),
    .A2(_07076_),
    .A3(_07098_),
    .B1(_07133_),
    .Y(_07208_));
 sky130_fd_sc_hd__mux2_1 _14534_ (.A0(\rbzero.wall_tracer.stepDistY[2] ),
    .A1(_07208_),
    .S(_07193_),
    .X(_07209_));
 sky130_fd_sc_hd__clkbuf_1 _14535_ (.A(_07209_),
    .X(_00420_));
 sky130_fd_sc_hd__or2_1 _14536_ (.A(_07133_),
    .B(_07052_),
    .X(_07210_));
 sky130_fd_sc_hd__nand2_1 _14537_ (.A(_07100_),
    .B(_07210_),
    .Y(_07211_));
 sky130_fd_sc_hd__mux2_1 _14538_ (.A0(\rbzero.wall_tracer.stepDistY[3] ),
    .A1(_07211_),
    .S(_07193_),
    .X(_07212_));
 sky130_fd_sc_hd__clkbuf_1 _14539_ (.A(_07212_),
    .X(_00421_));
 sky130_fd_sc_hd__buf_4 _14540_ (.A(_07099_),
    .X(_07213_));
 sky130_fd_sc_hd__nand2_1 _14541_ (.A(_05440_),
    .B(_07007_),
    .Y(_07214_));
 sky130_fd_sc_hd__a21oi_1 _14542_ (.A1(_07075_),
    .A2(_07088_),
    .B1(_07214_),
    .Y(_07215_));
 sky130_fd_sc_hd__a21oi_1 _14543_ (.A1(_07174_),
    .A2(_07092_),
    .B1(_07215_),
    .Y(_07216_));
 sky130_fd_sc_hd__nand2_1 _14544_ (.A(_07213_),
    .B(_07216_),
    .Y(_07217_));
 sky130_fd_sc_hd__mux2_1 _14545_ (.A0(\rbzero.wall_tracer.stepDistY[4] ),
    .A1(_07217_),
    .S(_07193_),
    .X(_07218_));
 sky130_fd_sc_hd__clkbuf_1 _14546_ (.A(_07218_),
    .X(_00422_));
 sky130_fd_sc_hd__nor2_1 _14547_ (.A(_05568_),
    .B(_07007_),
    .Y(_07219_));
 sky130_fd_sc_hd__o2bb2a_1 _14548_ (.A1_N(_07094_),
    .A2_N(_07219_),
    .B1(_07214_),
    .B2(_07085_),
    .X(_07220_));
 sky130_fd_sc_hd__nand2_1 _14549_ (.A(_07101_),
    .B(_07220_),
    .Y(_07221_));
 sky130_fd_sc_hd__mux2_1 _14550_ (.A0(\rbzero.wall_tracer.stepDistY[5] ),
    .A1(_07221_),
    .S(_07193_),
    .X(_07222_));
 sky130_fd_sc_hd__clkbuf_1 _14551_ (.A(_07222_),
    .X(_00423_));
 sky130_fd_sc_hd__nand3_1 _14552_ (.A(_06990_),
    .B(_06986_),
    .C(_06989_),
    .Y(_07223_));
 sky130_fd_sc_hd__or2_1 _14553_ (.A(_07082_),
    .B(_07214_),
    .X(_07224_));
 sky130_fd_sc_hd__o211ai_2 _14554_ (.A1(_07223_),
    .A2(_07096_),
    .B1(_07213_),
    .C1(_07224_),
    .Y(_07225_));
 sky130_fd_sc_hd__mux2_1 _14555_ (.A0(\rbzero.wall_tracer.stepDistY[6] ),
    .A1(_07225_),
    .S(_07193_),
    .X(_07226_));
 sky130_fd_sc_hd__clkbuf_1 _14556_ (.A(_07226_),
    .X(_00424_));
 sky130_fd_sc_hd__or4b_1 _14557_ (.A(_07029_),
    .B(_06985_),
    .C(_05568_),
    .D_N(_07031_),
    .X(_07227_));
 sky130_fd_sc_hd__a22o_1 _14558_ (.A1(_07007_),
    .A2(_07078_),
    .B1(_07214_),
    .B2(_07227_),
    .X(_07228_));
 sky130_fd_sc_hd__nand2_2 _14559_ (.A(_07101_),
    .B(_07228_),
    .Y(_07229_));
 sky130_fd_sc_hd__mux2_1 _14560_ (.A0(\rbzero.wall_tracer.stepDistY[7] ),
    .A1(_07229_),
    .S(_04925_),
    .X(_07230_));
 sky130_fd_sc_hd__clkbuf_1 _14561_ (.A(_07230_),
    .X(_00425_));
 sky130_fd_sc_hd__inv_2 _14562_ (.A(_07057_),
    .Y(_07231_));
 sky130_fd_sc_hd__a211o_1 _14563_ (.A1(_05401_),
    .A2(_06988_),
    .B1(_05406_),
    .C1(_06985_),
    .X(_07232_));
 sky130_fd_sc_hd__o211a_1 _14564_ (.A1(_05408_),
    .A2(_07231_),
    .B1(_07232_),
    .C1(_07075_),
    .X(_07233_));
 sky130_fd_sc_hd__a21oi_4 _14565_ (.A1(_07098_),
    .A2(_07233_),
    .B1(_07133_),
    .Y(_07234_));
 sky130_fd_sc_hd__mux2_1 _14566_ (.A0(\rbzero.wall_tracer.stepDistY[8] ),
    .A1(_07234_),
    .S(_04925_),
    .X(_07235_));
 sky130_fd_sc_hd__clkbuf_1 _14567_ (.A(_07235_),
    .X(_00426_));
 sky130_fd_sc_hd__inv_2 _14568_ (.A(_07213_),
    .Y(_07236_));
 sky130_fd_sc_hd__a31o_2 _14569_ (.A1(_05440_),
    .A2(_07007_),
    .A3(_07069_),
    .B1(_07236_),
    .X(_07237_));
 sky130_fd_sc_hd__mux2_1 _14570_ (.A0(\rbzero.wall_tracer.stepDistY[9] ),
    .A1(_07237_),
    .S(_04925_),
    .X(_07238_));
 sky130_fd_sc_hd__clkbuf_1 _14571_ (.A(_07238_),
    .X(_00427_));
 sky130_fd_sc_hd__nand2_1 _14572_ (.A(_06991_),
    .B(_07006_),
    .Y(_07239_));
 sky130_fd_sc_hd__or3_1 _14573_ (.A(_05416_),
    .B(_05408_),
    .C(_07239_),
    .X(_07240_));
 sky130_fd_sc_hd__nand2_1 _14574_ (.A(_07101_),
    .B(_07240_),
    .Y(_07241_));
 sky130_fd_sc_hd__mux2_1 _14575_ (.A0(\rbzero.wall_tracer.stepDistY[10] ),
    .A1(_07241_),
    .S(_04925_),
    .X(_07242_));
 sky130_fd_sc_hd__clkbuf_1 _14576_ (.A(_07242_),
    .X(_00428_));
 sky130_fd_sc_hd__and4_1 _14577_ (.A(_05440_),
    .B(_07007_),
    .C(_07038_),
    .D(_07101_),
    .X(_07243_));
 sky130_fd_sc_hd__mux2_1 _14578_ (.A0(\rbzero.wall_tracer.stepDistY[11] ),
    .A1(_07243_),
    .S(_04925_),
    .X(_07244_));
 sky130_fd_sc_hd__clkbuf_1 _14579_ (.A(_07244_),
    .X(_00429_));
 sky130_fd_sc_hd__buf_2 _14580_ (.A(_03799_),
    .X(_07245_));
 sky130_fd_sc_hd__clkbuf_4 _14581_ (.A(_05025_),
    .X(_07246_));
 sky130_fd_sc_hd__mux2_1 _14582_ (.A0(\rbzero.wall_tracer.trackDistX[-12] ),
    .A1(\rbzero.wall_tracer.trackDistY[-12] ),
    .S(_07246_),
    .X(_07247_));
 sky130_fd_sc_hd__and2_1 _14583_ (.A(_03797_),
    .B(_03778_),
    .X(_07248_));
 sky130_fd_sc_hd__clkbuf_4 _14584_ (.A(_07248_),
    .X(_07249_));
 sky130_fd_sc_hd__or2_1 _14585_ (.A(\rbzero.wall_tracer.visualWallDist[-12] ),
    .B(_07249_),
    .X(_07250_));
 sky130_fd_sc_hd__buf_2 _14586_ (.A(_03819_),
    .X(_07251_));
 sky130_fd_sc_hd__o211a_1 _14587_ (.A1(_07245_),
    .A2(_07247_),
    .B1(_07250_),
    .C1(_07251_),
    .X(_00430_));
 sky130_fd_sc_hd__buf_2 _14588_ (.A(_07248_),
    .X(_07252_));
 sky130_fd_sc_hd__clkbuf_4 _14589_ (.A(_07252_),
    .X(_07253_));
 sky130_fd_sc_hd__inv_2 _14590_ (.A(_05025_),
    .Y(_07254_));
 sky130_fd_sc_hd__nor2_1 _14591_ (.A(_05018_),
    .B(_07254_),
    .Y(_07255_));
 sky130_fd_sc_hd__o21ai_1 _14592_ (.A1(_04968_),
    .A2(_07246_),
    .B1(_07253_),
    .Y(_07256_));
 sky130_fd_sc_hd__clkbuf_4 _14593_ (.A(_03819_),
    .X(_07257_));
 sky130_fd_sc_hd__o221a_1 _14594_ (.A1(\rbzero.wall_tracer.visualWallDist[-11] ),
    .A2(_07253_),
    .B1(_07255_),
    .B2(_07256_),
    .C1(_07257_),
    .X(_00431_));
 sky130_fd_sc_hd__buf_4 _14595_ (.A(_05025_),
    .X(_07258_));
 sky130_fd_sc_hd__mux2_1 _14596_ (.A0(\rbzero.wall_tracer.trackDistX[-10] ),
    .A1(\rbzero.wall_tracer.trackDistY[-10] ),
    .S(_07258_),
    .X(_07259_));
 sky130_fd_sc_hd__clkinv_2 _14597_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .Y(_07260_));
 sky130_fd_sc_hd__nand2_1 _14598_ (.A(_07260_),
    .B(_03800_),
    .Y(_07261_));
 sky130_fd_sc_hd__o211a_1 _14599_ (.A1(_07245_),
    .A2(_07259_),
    .B1(_07261_),
    .C1(_07251_),
    .X(_00432_));
 sky130_fd_sc_hd__nor2_1 _14600_ (.A(_05020_),
    .B(_07254_),
    .Y(_07262_));
 sky130_fd_sc_hd__o21ai_1 _14601_ (.A1(_04965_),
    .A2(_07246_),
    .B1(_07249_),
    .Y(_07263_));
 sky130_fd_sc_hd__o221a_1 _14602_ (.A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A2(_07253_),
    .B1(_07262_),
    .B2(_07263_),
    .C1(_07257_),
    .X(_00433_));
 sky130_fd_sc_hd__nor2_1 _14603_ (.A(_05016_),
    .B(_07254_),
    .Y(_07264_));
 sky130_fd_sc_hd__o21ai_1 _14604_ (.A1(_04963_),
    .A2(_07246_),
    .B1(_07249_),
    .Y(_07265_));
 sky130_fd_sc_hd__clkbuf_4 _14605_ (.A(_03819_),
    .X(_07266_));
 sky130_fd_sc_hd__o221a_1 _14606_ (.A1(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A2(_07253_),
    .B1(_07264_),
    .B2(_07265_),
    .C1(_07266_),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _14607_ (.A0(\rbzero.wall_tracer.trackDistX[-7] ),
    .A1(\rbzero.wall_tracer.trackDistY[-7] ),
    .S(_07258_),
    .X(_07267_));
 sky130_fd_sc_hd__or2_1 _14608_ (.A(\rbzero.wall_tracer.visualWallDist[-7] ),
    .B(_07249_),
    .X(_07268_));
 sky130_fd_sc_hd__o211a_1 _14609_ (.A1(_07245_),
    .A2(_07267_),
    .B1(_07268_),
    .C1(_07251_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _14610_ (.A0(\rbzero.wall_tracer.trackDistX[-6] ),
    .A1(\rbzero.wall_tracer.trackDistY[-6] ),
    .S(_07258_),
    .X(_07269_));
 sky130_fd_sc_hd__or2_1 _14611_ (.A(\rbzero.wall_tracer.visualWallDist[-6] ),
    .B(_07249_),
    .X(_07270_));
 sky130_fd_sc_hd__o211a_1 _14612_ (.A1(_07245_),
    .A2(_07269_),
    .B1(_07270_),
    .C1(_07251_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _14613_ (.A0(\rbzero.wall_tracer.trackDistX[-5] ),
    .A1(\rbzero.wall_tracer.trackDistY[-5] ),
    .S(_07258_),
    .X(_07271_));
 sky130_fd_sc_hd__or2_1 _14614_ (.A(\rbzero.wall_tracer.visualWallDist[-5] ),
    .B(_07252_),
    .X(_07272_));
 sky130_fd_sc_hd__o211a_1 _14615_ (.A1(_07245_),
    .A2(_07271_),
    .B1(_07272_),
    .C1(_07251_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _14616_ (.A0(\rbzero.wall_tracer.trackDistX[-4] ),
    .A1(\rbzero.wall_tracer.trackDistY[-4] ),
    .S(_07258_),
    .X(_07273_));
 sky130_fd_sc_hd__or2_1 _14617_ (.A(\rbzero.wall_tracer.visualWallDist[-4] ),
    .B(_07252_),
    .X(_07274_));
 sky130_fd_sc_hd__o211a_1 _14618_ (.A1(_07245_),
    .A2(_07273_),
    .B1(_07274_),
    .C1(_07251_),
    .X(_00438_));
 sky130_fd_sc_hd__inv_2 _14619_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .Y(_07275_));
 sky130_fd_sc_hd__nor2_1 _14620_ (.A(_07275_),
    .B(_07254_),
    .Y(_07276_));
 sky130_fd_sc_hd__o21ai_1 _14621_ (.A1(_04947_),
    .A2(_07246_),
    .B1(_07249_),
    .Y(_07277_));
 sky130_fd_sc_hd__o221a_1 _14622_ (.A1(\rbzero.wall_tracer.visualWallDist[-3] ),
    .A2(_07253_),
    .B1(_07276_),
    .B2(_07277_),
    .C1(_07266_),
    .X(_00439_));
 sky130_fd_sc_hd__nor2_1 _14623_ (.A(_04954_),
    .B(_07254_),
    .Y(_07278_));
 sky130_fd_sc_hd__o21ai_1 _14624_ (.A1(_04950_),
    .A2(_07246_),
    .B1(_07249_),
    .Y(_07279_));
 sky130_fd_sc_hd__o221a_1 _14625_ (.A1(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A2(_07253_),
    .B1(_07278_),
    .B2(_07279_),
    .C1(_07266_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _14626_ (.A0(\rbzero.wall_tracer.trackDistX[-1] ),
    .A1(\rbzero.wall_tracer.trackDistY[-1] ),
    .S(_07258_),
    .X(_07280_));
 sky130_fd_sc_hd__or2_1 _14627_ (.A(\rbzero.wall_tracer.visualWallDist[-1] ),
    .B(_07252_),
    .X(_07281_));
 sky130_fd_sc_hd__o211a_1 _14628_ (.A1(_07245_),
    .A2(_07280_),
    .B1(_07281_),
    .C1(_07251_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _14629_ (.A0(\rbzero.wall_tracer.trackDistX[0] ),
    .A1(\rbzero.wall_tracer.trackDistY[0] ),
    .S(_07258_),
    .X(_07282_));
 sky130_fd_sc_hd__or2_1 _14630_ (.A(\rbzero.wall_tracer.visualWallDist[0] ),
    .B(_07252_),
    .X(_07283_));
 sky130_fd_sc_hd__o211a_1 _14631_ (.A1(_07245_),
    .A2(_07282_),
    .B1(_07283_),
    .C1(_07251_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _14632_ (.A0(\rbzero.wall_tracer.trackDistX[1] ),
    .A1(\rbzero.wall_tracer.trackDistY[1] ),
    .S(_07258_),
    .X(_07284_));
 sky130_fd_sc_hd__or2_1 _14633_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_07252_),
    .X(_07285_));
 sky130_fd_sc_hd__o211a_1 _14634_ (.A1(_07245_),
    .A2(_07284_),
    .B1(_07285_),
    .C1(_07251_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _14635_ (.A0(\rbzero.wall_tracer.trackDistX[2] ),
    .A1(\rbzero.wall_tracer.trackDistY[2] ),
    .S(_07258_),
    .X(_07286_));
 sky130_fd_sc_hd__or2_1 _14636_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_07252_),
    .X(_07287_));
 sky130_fd_sc_hd__o211a_1 _14637_ (.A1(_07245_),
    .A2(_07286_),
    .B1(_07287_),
    .C1(_07251_),
    .X(_00444_));
 sky130_fd_sc_hd__nor2_1 _14638_ (.A(_04941_),
    .B(_07254_),
    .Y(_07288_));
 sky130_fd_sc_hd__o21ai_1 _14639_ (.A1(_04985_),
    .A2(_07246_),
    .B1(_07249_),
    .Y(_07289_));
 sky130_fd_sc_hd__o221a_1 _14640_ (.A1(\rbzero.wall_tracer.visualWallDist[3] ),
    .A2(_07253_),
    .B1(_07288_),
    .B2(_07289_),
    .C1(_07266_),
    .X(_00445_));
 sky130_fd_sc_hd__nor2_1 _14641_ (.A(_05001_),
    .B(_07254_),
    .Y(_07290_));
 sky130_fd_sc_hd__inv_2 _14642_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .Y(_07291_));
 sky130_fd_sc_hd__o21ai_1 _14643_ (.A1(_07291_),
    .A2(_07246_),
    .B1(_07249_),
    .Y(_07292_));
 sky130_fd_sc_hd__o221a_1 _14644_ (.A1(\rbzero.wall_tracer.visualWallDist[4] ),
    .A2(_07253_),
    .B1(_07290_),
    .B2(_07292_),
    .C1(_07266_),
    .X(_00446_));
 sky130_fd_sc_hd__nor2_1 _14645_ (.A(_05002_),
    .B(_07254_),
    .Y(_07293_));
 sky130_fd_sc_hd__inv_2 _14646_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .Y(_07294_));
 sky130_fd_sc_hd__o21ai_1 _14647_ (.A1(_07294_),
    .A2(_07246_),
    .B1(_07249_),
    .Y(_07295_));
 sky130_fd_sc_hd__o221a_1 _14648_ (.A1(\rbzero.wall_tracer.visualWallDist[5] ),
    .A2(_07253_),
    .B1(_07293_),
    .B2(_07295_),
    .C1(_07266_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _14649_ (.A0(\rbzero.wall_tracer.trackDistX[6] ),
    .A1(\rbzero.wall_tracer.trackDistY[6] ),
    .S(_07258_),
    .X(_07296_));
 sky130_fd_sc_hd__or2_1 _14650_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_07252_),
    .X(_07297_));
 sky130_fd_sc_hd__o211a_1 _14651_ (.A1(_03800_),
    .A2(_07296_),
    .B1(_07297_),
    .C1(_07257_),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _14652_ (.A0(\rbzero.wall_tracer.trackDistX[7] ),
    .A1(\rbzero.wall_tracer.trackDistY[7] ),
    .S(_05025_),
    .X(_07298_));
 sky130_fd_sc_hd__or2_1 _14653_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_07252_),
    .X(_07299_));
 sky130_fd_sc_hd__o211a_1 _14654_ (.A1(_03800_),
    .A2(_07298_),
    .B1(_07299_),
    .C1(_07257_),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _14655_ (.A0(\rbzero.wall_tracer.trackDistX[8] ),
    .A1(\rbzero.wall_tracer.trackDistY[8] ),
    .S(_05025_),
    .X(_07300_));
 sky130_fd_sc_hd__nand2_1 _14656_ (.A(_05290_),
    .B(_03800_),
    .Y(_07301_));
 sky130_fd_sc_hd__o211a_1 _14657_ (.A1(_03800_),
    .A2(_07300_),
    .B1(_07301_),
    .C1(_07257_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _14658_ (.A0(\rbzero.wall_tracer.trackDistX[9] ),
    .A1(\rbzero.wall_tracer.trackDistY[9] ),
    .S(_05025_),
    .X(_07302_));
 sky130_fd_sc_hd__or2_1 _14659_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_07252_),
    .X(_07303_));
 sky130_fd_sc_hd__o211a_1 _14660_ (.A1(_03800_),
    .A2(_07302_),
    .B1(_07303_),
    .C1(_07257_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _14661_ (.A0(\rbzero.wall_tracer.trackDistX[10] ),
    .A1(\rbzero.wall_tracer.trackDistY[10] ),
    .S(_05025_),
    .X(_07304_));
 sky130_fd_sc_hd__nand2_1 _14662_ (.A(_05301_),
    .B(_03800_),
    .Y(_07305_));
 sky130_fd_sc_hd__o211a_1 _14663_ (.A1(_03800_),
    .A2(_07304_),
    .B1(_07305_),
    .C1(_07257_),
    .X(_00452_));
 sky130_fd_sc_hd__a21o_1 _14664_ (.A1(\rbzero.wall_tracer.trackDistY[11] ),
    .A2(\rbzero.wall_tracer.trackDistX[11] ),
    .B1(_03799_),
    .X(_07306_));
 sky130_fd_sc_hd__o211a_1 _14665_ (.A1(\rbzero.wall_tracer.visualWallDist[11] ),
    .A2(_07253_),
    .B1(_07306_),
    .C1(_07257_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _14666_ (.A0(\rbzero.wall_tracer.stepDistX[-12] ),
    .A1(_07118_),
    .S(_00008_),
    .X(_07307_));
 sky130_fd_sc_hd__clkbuf_1 _14667_ (.A(_07307_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _14668_ (.A0(\rbzero.wall_tracer.stepDistX[-11] ),
    .A1(_07136_),
    .S(_00008_),
    .X(_07308_));
 sky130_fd_sc_hd__clkbuf_1 _14669_ (.A(_07308_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _14670_ (.A0(\rbzero.wall_tracer.stepDistX[-10] ),
    .A1(_07147_),
    .S(_00008_),
    .X(_07309_));
 sky130_fd_sc_hd__clkbuf_1 _14671_ (.A(_07309_),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _14672_ (.A0(\rbzero.wall_tracer.stepDistX[-9] ),
    .A1(_07157_),
    .S(_00008_),
    .X(_07310_));
 sky130_fd_sc_hd__clkbuf_1 _14673_ (.A(_07310_),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _14674_ (.A0(\rbzero.wall_tracer.stepDistX[-8] ),
    .A1(_07165_),
    .S(_00008_),
    .X(_07311_));
 sky130_fd_sc_hd__clkbuf_1 _14675_ (.A(_07311_),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _14676_ (.A0(\rbzero.wall_tracer.stepDistX[-7] ),
    .A1(_07172_),
    .S(_00008_),
    .X(_07312_));
 sky130_fd_sc_hd__clkbuf_1 _14677_ (.A(_07312_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _14678_ (.A0(\rbzero.wall_tracer.stepDistX[-6] ),
    .A1(_07180_),
    .S(_00008_),
    .X(_07313_));
 sky130_fd_sc_hd__clkbuf_1 _14679_ (.A(_07313_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _14680_ (.A0(\rbzero.wall_tracer.stepDistX[-5] ),
    .A1(_07185_),
    .S(_00008_),
    .X(_07314_));
 sky130_fd_sc_hd__clkbuf_1 _14681_ (.A(_07314_),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _14682_ (.A0(\rbzero.wall_tracer.stepDistX[-4] ),
    .A1(_07189_),
    .S(_00008_),
    .X(_07315_));
 sky130_fd_sc_hd__clkbuf_1 _14683_ (.A(_07315_),
    .X(_00462_));
 sky130_fd_sc_hd__buf_4 _14684_ (.A(_04931_),
    .X(_07316_));
 sky130_fd_sc_hd__mux2_1 _14685_ (.A0(\rbzero.wall_tracer.stepDistX[-3] ),
    .A1(_07192_),
    .S(_07316_),
    .X(_07317_));
 sky130_fd_sc_hd__clkbuf_1 _14686_ (.A(_07317_),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _14687_ (.A0(\rbzero.wall_tracer.stepDistX[-2] ),
    .A1(_07196_),
    .S(_07316_),
    .X(_07318_));
 sky130_fd_sc_hd__clkbuf_1 _14688_ (.A(_07318_),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _14689_ (.A0(\rbzero.wall_tracer.stepDistX[-1] ),
    .A1(_07199_),
    .S(_07316_),
    .X(_07319_));
 sky130_fd_sc_hd__clkbuf_1 _14690_ (.A(_07319_),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _14691_ (.A0(\rbzero.wall_tracer.stepDistX[0] ),
    .A1(_07202_),
    .S(_07316_),
    .X(_07320_));
 sky130_fd_sc_hd__clkbuf_1 _14692_ (.A(_07320_),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _14693_ (.A0(\rbzero.wall_tracer.stepDistX[1] ),
    .A1(_07206_),
    .S(_07316_),
    .X(_07321_));
 sky130_fd_sc_hd__clkbuf_1 _14694_ (.A(_07321_),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _14695_ (.A0(\rbzero.wall_tracer.stepDistX[2] ),
    .A1(_07208_),
    .S(_07316_),
    .X(_07322_));
 sky130_fd_sc_hd__clkbuf_1 _14696_ (.A(_07322_),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _14697_ (.A0(\rbzero.wall_tracer.stepDistX[3] ),
    .A1(_07211_),
    .S(_07316_),
    .X(_07323_));
 sky130_fd_sc_hd__clkbuf_1 _14698_ (.A(_07323_),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _14699_ (.A0(\rbzero.wall_tracer.stepDistX[4] ),
    .A1(_07217_),
    .S(_07316_),
    .X(_07324_));
 sky130_fd_sc_hd__clkbuf_1 _14700_ (.A(_07324_),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _14701_ (.A0(\rbzero.wall_tracer.stepDistX[5] ),
    .A1(_07221_),
    .S(_07316_),
    .X(_07325_));
 sky130_fd_sc_hd__clkbuf_1 _14702_ (.A(_07325_),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _14703_ (.A0(\rbzero.wall_tracer.stepDistX[6] ),
    .A1(_07225_),
    .S(_07316_),
    .X(_07326_));
 sky130_fd_sc_hd__clkbuf_1 _14704_ (.A(_07326_),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _14705_ (.A0(\rbzero.wall_tracer.stepDistX[7] ),
    .A1(_07229_),
    .S(_04931_),
    .X(_07327_));
 sky130_fd_sc_hd__clkbuf_1 _14706_ (.A(_07327_),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _14707_ (.A0(\rbzero.wall_tracer.stepDistX[8] ),
    .A1(_07234_),
    .S(_04931_),
    .X(_07328_));
 sky130_fd_sc_hd__clkbuf_1 _14708_ (.A(_07328_),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _14709_ (.A0(\rbzero.wall_tracer.stepDistX[9] ),
    .A1(_07237_),
    .S(_04931_),
    .X(_07329_));
 sky130_fd_sc_hd__clkbuf_1 _14710_ (.A(_07329_),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _14711_ (.A0(\rbzero.wall_tracer.stepDistX[10] ),
    .A1(_07241_),
    .S(_04931_),
    .X(_07330_));
 sky130_fd_sc_hd__clkbuf_1 _14712_ (.A(_07330_),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _14713_ (.A0(\rbzero.wall_tracer.stepDistX[11] ),
    .A1(_07243_),
    .S(_04931_),
    .X(_07331_));
 sky130_fd_sc_hd__clkbuf_1 _14714_ (.A(_07331_),
    .X(_00477_));
 sky130_fd_sc_hd__buf_4 _14715_ (.A(_04940_),
    .X(_07332_));
 sky130_fd_sc_hd__nor2_1 _14716_ (.A(_07332_),
    .B(_03777_),
    .Y(_07333_));
 sky130_fd_sc_hd__a32o_1 _14717_ (.A1(_03819_),
    .A2(_03756_),
    .A3(_07333_),
    .B1(_05026_),
    .B2(\rbzero.wall_tracer.wall[0] ),
    .X(_00478_));
 sky130_fd_sc_hd__a32o_1 _14718_ (.A1(_03819_),
    .A2(_03764_),
    .A3(_07333_),
    .B1(_05026_),
    .B2(\rbzero.wall_tracer.wall[1] ),
    .X(_00479_));
 sky130_fd_sc_hd__inv_2 _14719_ (.A(\rbzero.wall_tracer.side ),
    .Y(_07334_));
 sky130_fd_sc_hd__nand2_1 _14720_ (.A(_07334_),
    .B(_03799_),
    .Y(_07335_));
 sky130_fd_sc_hd__o211a_1 _14721_ (.A1(_03800_),
    .A2(_07246_),
    .B1(_07335_),
    .C1(_07257_),
    .X(_00480_));
 sky130_fd_sc_hd__buf_4 _14722_ (.A(\rbzero.wall_tracer.state[3] ),
    .X(_07336_));
 sky130_fd_sc_hd__buf_4 _14723_ (.A(_07336_),
    .X(_07337_));
 sky130_fd_sc_hd__buf_4 _14724_ (.A(_07337_),
    .X(_07338_));
 sky130_fd_sc_hd__inv_2 _14725_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .Y(_07339_));
 sky130_fd_sc_hd__inv_2 _14726_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .Y(_07340_));
 sky130_fd_sc_hd__buf_2 _14727_ (.A(\rbzero.wall_tracer.side ),
    .X(_07341_));
 sky130_fd_sc_hd__buf_2 _14728_ (.A(_07341_),
    .X(_07342_));
 sky130_fd_sc_hd__clkbuf_4 _14729_ (.A(_07342_),
    .X(_07343_));
 sky130_fd_sc_hd__mux2_1 _14730_ (.A0(_07339_),
    .A1(_07340_),
    .S(_07343_),
    .X(_07344_));
 sky130_fd_sc_hd__a31o_1 _14731_ (.A1(_07100_),
    .A2(_07187_),
    .A3(_07188_),
    .B1(_07336_),
    .X(_07345_));
 sky130_fd_sc_hd__buf_2 _14732_ (.A(\rbzero.wall_tracer.state[3] ),
    .X(_07346_));
 sky130_fd_sc_hd__mux2_1 _14733_ (.A0(_05085_),
    .A1(_05226_),
    .S(_07341_),
    .X(_07347_));
 sky130_fd_sc_hd__nand2_1 _14734_ (.A(_07346_),
    .B(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__clkbuf_4 _14735_ (.A(\rbzero.wall_tracer.state[13] ),
    .X(_07349_));
 sky130_fd_sc_hd__a21o_1 _14736_ (.A1(_07345_),
    .A2(_07348_),
    .B1(_07349_),
    .X(_07350_));
 sky130_fd_sc_hd__clkbuf_4 _14737_ (.A(\rbzero.wall_tracer.state[13] ),
    .X(_07351_));
 sky130_fd_sc_hd__buf_4 _14738_ (.A(\rbzero.wall_tracer.state[6] ),
    .X(_07352_));
 sky130_fd_sc_hd__a21oi_2 _14739_ (.A1(_07351_),
    .A2(\rbzero.wall_tracer.stepDistY[-4] ),
    .B1(_07352_),
    .Y(_07353_));
 sky130_fd_sc_hd__nor2_1 _14740_ (.A(_04927_),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .Y(_07354_));
 sky130_fd_sc_hd__a21o_2 _14741_ (.A1(_07350_),
    .A2(_07353_),
    .B1(_07354_),
    .X(_07355_));
 sky130_fd_sc_hd__buf_4 _14742_ (.A(_07352_),
    .X(_07356_));
 sky130_fd_sc_hd__or3_1 _14743_ (.A(\rbzero.debug_overlay.playerY[-7] ),
    .B(\rbzero.debug_overlay.playerY[-8] ),
    .C(\rbzero.debug_overlay.playerY[-9] ),
    .X(_07357_));
 sky130_fd_sc_hd__or2_1 _14744_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_07357_),
    .X(_07358_));
 sky130_fd_sc_hd__nand2_1 _14745_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_07357_),
    .Y(_07359_));
 sky130_fd_sc_hd__and2_1 _14746_ (.A(_07358_),
    .B(_07359_),
    .X(_07360_));
 sky130_fd_sc_hd__nand2_1 _14747_ (.A(_07339_),
    .B(_05113_),
    .Y(_07361_));
 sky130_fd_sc_hd__o211a_1 _14748_ (.A1(_05113_),
    .A2(_07360_),
    .B1(_07361_),
    .C1(_07351_),
    .X(_07362_));
 sky130_fd_sc_hd__and2_1 _14749_ (.A(\rbzero.wall_tracer.visualWallDist[-6] ),
    .B(_03793_),
    .X(_07363_));
 sky130_fd_sc_hd__or3_1 _14750_ (.A(\rbzero.debug_overlay.playerX[-7] ),
    .B(\rbzero.debug_overlay.playerX[-8] ),
    .C(\rbzero.debug_overlay.playerX[-9] ),
    .X(_07364_));
 sky130_fd_sc_hd__or2_1 _14751_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .B(_07364_),
    .X(_07365_));
 sky130_fd_sc_hd__nand2_1 _14752_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .B(_07364_),
    .Y(_07366_));
 sky130_fd_sc_hd__nand2_1 _14753_ (.A(_07365_),
    .B(_07366_),
    .Y(_07367_));
 sky130_fd_sc_hd__inv_2 _14754_ (.A(_05273_),
    .Y(_07368_));
 sky130_fd_sc_hd__or4_1 _14755_ (.A(\rbzero.wall_tracer.rayAddendX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .C(\rbzero.wall_tracer.rayAddendX[-2] ),
    .D(_05258_),
    .X(_07369_));
 sky130_fd_sc_hd__or4_1 _14756_ (.A(_05236_),
    .B(_05247_),
    .C(_05242_),
    .D(_07369_),
    .X(_07370_));
 sky130_fd_sc_hd__or4b_1 _14757_ (.A(_05226_),
    .B(_07370_),
    .C(_05221_),
    .D_N(_05230_),
    .X(_07371_));
 sky130_fd_sc_hd__or3b_1 _14758_ (.A(_07371_),
    .B(_05267_),
    .C_N(_05215_),
    .X(_07372_));
 sky130_fd_sc_hd__and3b_1 _14759_ (.A_N(_07372_),
    .B(_05203_),
    .C(_05210_),
    .X(_07373_));
 sky130_fd_sc_hd__a31oi_4 _14760_ (.A1(_05196_),
    .A2(_07368_),
    .A3(_07373_),
    .B1(_05186_),
    .Y(_07374_));
 sky130_fd_sc_hd__mux2_1 _14761_ (.A0(_07340_),
    .A1(_07367_),
    .S(_07374_),
    .X(_07375_));
 sky130_fd_sc_hd__nand2_1 _14762_ (.A(_04935_),
    .B(_07375_),
    .Y(_07376_));
 sky130_fd_sc_hd__o31ai_4 _14763_ (.A1(_07356_),
    .A2(_07362_),
    .A3(_07363_),
    .B1(_07376_),
    .Y(_07377_));
 sky130_fd_sc_hd__buf_2 _14764_ (.A(_07377_),
    .X(_07378_));
 sky130_fd_sc_hd__clkbuf_4 _14765_ (.A(_07378_),
    .X(_07379_));
 sky130_fd_sc_hd__nor2_1 _14766_ (.A(_07355_),
    .B(_07379_),
    .Y(_07380_));
 sky130_fd_sc_hd__a21o_1 _14767_ (.A1(_07213_),
    .A2(_07184_),
    .B1(_07336_),
    .X(_07381_));
 sky130_fd_sc_hd__nor2_1 _14768_ (.A(_07341_),
    .B(_05091_),
    .Y(_07382_));
 sky130_fd_sc_hd__a211o_1 _14769_ (.A1(_07341_),
    .A2(_05230_),
    .B1(_07382_),
    .C1(_04932_),
    .X(_07383_));
 sky130_fd_sc_hd__a21o_1 _14770_ (.A1(_07381_),
    .A2(_07383_),
    .B1(_07349_),
    .X(_07384_));
 sky130_fd_sc_hd__a21oi_2 _14771_ (.A1(_07351_),
    .A2(\rbzero.wall_tracer.stepDistY[-5] ),
    .B1(_07352_),
    .Y(_07385_));
 sky130_fd_sc_hd__nor2_1 _14772_ (.A(_04927_),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .Y(_07386_));
 sky130_fd_sc_hd__a21o_2 _14773_ (.A1(_07384_),
    .A2(_07385_),
    .B1(_07386_),
    .X(_07387_));
 sky130_fd_sc_hd__buf_2 _14774_ (.A(_07387_),
    .X(_07388_));
 sky130_fd_sc_hd__inv_2 _14775_ (.A(\rbzero.debug_overlay.playerY[-5] ),
    .Y(_07389_));
 sky130_fd_sc_hd__xnor2_1 _14776_ (.A(_07389_),
    .B(_07358_),
    .Y(_07390_));
 sky130_fd_sc_hd__nand2_1 _14777_ (.A(_07389_),
    .B(_05113_),
    .Y(_07391_));
 sky130_fd_sc_hd__o211a_1 _14778_ (.A1(_05113_),
    .A2(_07390_),
    .B1(_07391_),
    .C1(_07351_),
    .X(_07392_));
 sky130_fd_sc_hd__and2_1 _14779_ (.A(\rbzero.wall_tracer.visualWallDist[-5] ),
    .B(_03793_),
    .X(_07393_));
 sky130_fd_sc_hd__inv_2 _14780_ (.A(\rbzero.debug_overlay.playerX[-5] ),
    .Y(_07394_));
 sky130_fd_sc_hd__xnor2_1 _14781_ (.A(\rbzero.debug_overlay.playerX[-5] ),
    .B(_07365_),
    .Y(_07395_));
 sky130_fd_sc_hd__mux2_1 _14782_ (.A0(_07394_),
    .A1(_07395_),
    .S(_07374_),
    .X(_07396_));
 sky130_fd_sc_hd__nand2_1 _14783_ (.A(_04935_),
    .B(_07396_),
    .Y(_07397_));
 sky130_fd_sc_hd__o31ai_4 _14784_ (.A1(_07356_),
    .A2(_07392_),
    .A3(_07393_),
    .B1(_07397_),
    .Y(_07398_));
 sky130_fd_sc_hd__clkbuf_4 _14785_ (.A(_07398_),
    .X(_07399_));
 sky130_fd_sc_hd__buf_4 _14786_ (.A(_07399_),
    .X(_07400_));
 sky130_fd_sc_hd__nor2_1 _14787_ (.A(_07388_),
    .B(_07400_),
    .Y(_07401_));
 sky130_fd_sc_hd__or4_1 _14788_ (.A(_07355_),
    .B(_07378_),
    .C(_07387_),
    .D(_07399_),
    .X(_07402_));
 sky130_fd_sc_hd__o21ai_1 _14789_ (.A1(_07380_),
    .A2(_07401_),
    .B1(_07402_),
    .Y(_07403_));
 sky130_fd_sc_hd__or3_1 _14790_ (.A(\rbzero.debug_overlay.playerY[-4] ),
    .B(\rbzero.debug_overlay.playerY[-5] ),
    .C(_07358_),
    .X(_07404_));
 sky130_fd_sc_hd__o21ai_1 _14791_ (.A1(\rbzero.debug_overlay.playerY[-5] ),
    .A2(_07358_),
    .B1(\rbzero.debug_overlay.playerY[-4] ),
    .Y(_07405_));
 sky130_fd_sc_hd__and2_1 _14792_ (.A(_07404_),
    .B(_07405_),
    .X(_07406_));
 sky130_fd_sc_hd__mux2_1 _14793_ (.A0(_07406_),
    .A1(\rbzero.debug_overlay.playerY[-4] ),
    .S(_05113_),
    .X(_07407_));
 sky130_fd_sc_hd__clkbuf_4 _14794_ (.A(_07349_),
    .X(_07408_));
 sky130_fd_sc_hd__mux2_1 _14795_ (.A0(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A1(_07407_),
    .S(_07408_),
    .X(_07409_));
 sky130_fd_sc_hd__inv_2 _14796_ (.A(\rbzero.debug_overlay.playerX[-4] ),
    .Y(_07410_));
 sky130_fd_sc_hd__or3_1 _14797_ (.A(\rbzero.debug_overlay.playerX[-4] ),
    .B(\rbzero.debug_overlay.playerX[-5] ),
    .C(_07365_),
    .X(_07411_));
 sky130_fd_sc_hd__o21ai_1 _14798_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_07365_),
    .B1(\rbzero.debug_overlay.playerX[-4] ),
    .Y(_07412_));
 sky130_fd_sc_hd__nand2_1 _14799_ (.A(_07411_),
    .B(_07412_),
    .Y(_07413_));
 sky130_fd_sc_hd__mux2_1 _14800_ (.A0(_07410_),
    .A1(_07413_),
    .S(_07374_),
    .X(_07414_));
 sky130_fd_sc_hd__nand2_1 _14801_ (.A(_04936_),
    .B(_07414_),
    .Y(_07415_));
 sky130_fd_sc_hd__o21ai_4 _14802_ (.A1(_04936_),
    .A2(_07409_),
    .B1(_07415_),
    .Y(_07416_));
 sky130_fd_sc_hd__a21o_1 _14803_ (.A1(_07213_),
    .A2(_07179_),
    .B1(_07346_),
    .X(_07417_));
 sky130_fd_sc_hd__mux2_1 _14804_ (.A0(_05089_),
    .A1(_05236_),
    .S(_07341_),
    .X(_07418_));
 sky130_fd_sc_hd__nand2_1 _14805_ (.A(_07346_),
    .B(_07418_),
    .Y(_07419_));
 sky130_fd_sc_hd__a21o_1 _14806_ (.A1(_07417_),
    .A2(_07419_),
    .B1(_07349_),
    .X(_07420_));
 sky130_fd_sc_hd__a21oi_2 _14807_ (.A1(_07351_),
    .A2(\rbzero.wall_tracer.stepDistY[-6] ),
    .B1(_07352_),
    .Y(_07421_));
 sky130_fd_sc_hd__nor2_1 _14808_ (.A(_04927_),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .Y(_07422_));
 sky130_fd_sc_hd__a21o_1 _14809_ (.A1(_07420_),
    .A2(_07421_),
    .B1(_07422_),
    .X(_07423_));
 sky130_fd_sc_hd__buf_2 _14810_ (.A(_07423_),
    .X(_07424_));
 sky130_fd_sc_hd__or2_1 _14811_ (.A(_07416_),
    .B(_07424_),
    .X(_07425_));
 sky130_fd_sc_hd__xnor2_1 _14812_ (.A(_07403_),
    .B(_07425_),
    .Y(_07426_));
 sky130_fd_sc_hd__xor2_1 _14813_ (.A(\rbzero.debug_overlay.playerY[-8] ),
    .B(\rbzero.debug_overlay.playerY[-9] ),
    .X(_07427_));
 sky130_fd_sc_hd__mux2_1 _14814_ (.A0(_07427_),
    .A1(\rbzero.debug_overlay.playerY[-8] ),
    .S(_05113_),
    .X(_07428_));
 sky130_fd_sc_hd__nand2_1 _14815_ (.A(_07349_),
    .B(_07428_),
    .Y(_07429_));
 sky130_fd_sc_hd__a21oi_1 _14816_ (.A1(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A2(_03793_),
    .B1(\rbzero.wall_tracer.state[6] ),
    .Y(_07430_));
 sky130_fd_sc_hd__inv_2 _14817_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .Y(_07431_));
 sky130_fd_sc_hd__xnor2_1 _14818_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .B(\rbzero.debug_overlay.playerX[-9] ),
    .Y(_07432_));
 sky130_fd_sc_hd__mux2_1 _14819_ (.A0(_07431_),
    .A1(_07432_),
    .S(_07374_),
    .X(_07433_));
 sky130_fd_sc_hd__a22o_1 _14820_ (.A1(_07429_),
    .A2(_07430_),
    .B1(_07433_),
    .B2(_07352_),
    .X(_07434_));
 sky130_fd_sc_hd__buf_2 _14821_ (.A(_07434_),
    .X(_07435_));
 sky130_fd_sc_hd__a21o_1 _14822_ (.A1(_07100_),
    .A2(_07191_),
    .B1(_07336_),
    .X(_07436_));
 sky130_fd_sc_hd__mux2_1 _14823_ (.A0(_05084_),
    .A1(_05221_),
    .S(\rbzero.wall_tracer.side ),
    .X(_07437_));
 sky130_fd_sc_hd__nand2_1 _14824_ (.A(_07336_),
    .B(_07437_),
    .Y(_07438_));
 sky130_fd_sc_hd__a21o_1 _14825_ (.A1(_07436_),
    .A2(_07438_),
    .B1(\rbzero.wall_tracer.state[13] ),
    .X(_07439_));
 sky130_fd_sc_hd__a21oi_2 _14826_ (.A1(\rbzero.wall_tracer.state[13] ),
    .A2(\rbzero.wall_tracer.stepDistY[-3] ),
    .B1(\rbzero.wall_tracer.state[6] ),
    .Y(_07440_));
 sky130_fd_sc_hd__nor2_1 _14827_ (.A(_04927_),
    .B(\rbzero.wall_tracer.stepDistX[-3] ),
    .Y(_07441_));
 sky130_fd_sc_hd__a21o_1 _14828_ (.A1(_07439_),
    .A2(_07440_),
    .B1(_07441_),
    .X(_07442_));
 sky130_fd_sc_hd__nand2_2 _14829_ (.A(\rbzero.wall_tracer.visualWallDist[-12] ),
    .B(_03795_),
    .Y(_07443_));
 sky130_fd_sc_hd__nand3_1 _14830_ (.A(_07099_),
    .B(_07195_),
    .C(_07198_),
    .Y(_07444_));
 sky130_fd_sc_hd__a21o_2 _14831_ (.A1(_07202_),
    .A2(_07444_),
    .B1(_07206_),
    .X(_07445_));
 sky130_fd_sc_hd__o211a_1 _14832_ (.A1(_07177_),
    .A2(_07162_),
    .B1(_07201_),
    .C1(_07100_),
    .X(_07446_));
 sky130_fd_sc_hd__and3_1 _14833_ (.A(_07100_),
    .B(_07204_),
    .C(_07205_),
    .X(_07447_));
 sky130_fd_sc_hd__and3_1 _14834_ (.A(_07099_),
    .B(_07195_),
    .C(_07198_),
    .X(_07448_));
 sky130_fd_sc_hd__or3_1 _14835_ (.A(_07446_),
    .B(_07447_),
    .C(_07448_),
    .X(_07449_));
 sky130_fd_sc_hd__a21oi_2 _14836_ (.A1(_07445_),
    .A2(_07449_),
    .B1(_07337_),
    .Y(_07450_));
 sky130_fd_sc_hd__nand2_1 _14837_ (.A(_07342_),
    .B(_05203_),
    .Y(_07451_));
 sky130_fd_sc_hd__or2_1 _14838_ (.A(_07342_),
    .B(_05080_),
    .X(_07452_));
 sky130_fd_sc_hd__buf_4 _14839_ (.A(_07351_),
    .X(_07453_));
 sky130_fd_sc_hd__a31o_1 _14840_ (.A1(_07337_),
    .A2(_07451_),
    .A3(_07452_),
    .B1(_07453_),
    .X(_07454_));
 sky130_fd_sc_hd__o221ai_4 _14841_ (.A1(_03795_),
    .A2(\rbzero.wall_tracer.stepDistY[1] ),
    .B1(_07450_),
    .B2(_07454_),
    .C1(_04928_),
    .Y(_07455_));
 sky130_fd_sc_hd__or4_1 _14842_ (.A(_07435_),
    .B(_07442_),
    .C(_07443_),
    .D(_07455_),
    .X(_07456_));
 sky130_fd_sc_hd__o21ai_1 _14843_ (.A1(\rbzero.debug_overlay.playerY[-8] ),
    .A2(\rbzero.debug_overlay.playerY[-9] ),
    .B1(\rbzero.debug_overlay.playerY[-7] ),
    .Y(_07457_));
 sky130_fd_sc_hd__and2_1 _14844_ (.A(_07357_),
    .B(_07457_),
    .X(_07458_));
 sky130_fd_sc_hd__mux2_1 _14845_ (.A0(_07458_),
    .A1(\rbzero.debug_overlay.playerY[-7] ),
    .S(_05113_),
    .X(_07459_));
 sky130_fd_sc_hd__nand2_1 _14846_ (.A(_07453_),
    .B(_07459_),
    .Y(_07460_));
 sky130_fd_sc_hd__a21oi_1 _14847_ (.A1(\rbzero.wall_tracer.visualWallDist[-7] ),
    .A2(_03795_),
    .B1(_04936_),
    .Y(_07461_));
 sky130_fd_sc_hd__inv_2 _14848_ (.A(\rbzero.debug_overlay.playerX[-7] ),
    .Y(_07462_));
 sky130_fd_sc_hd__o21ai_1 _14849_ (.A1(\rbzero.debug_overlay.playerX[-8] ),
    .A2(\rbzero.debug_overlay.playerX[-9] ),
    .B1(\rbzero.debug_overlay.playerX[-7] ),
    .Y(_07463_));
 sky130_fd_sc_hd__nand2_1 _14850_ (.A(_07364_),
    .B(_07463_),
    .Y(_07464_));
 sky130_fd_sc_hd__mux2_1 _14851_ (.A0(_07462_),
    .A1(_07464_),
    .S(_07374_),
    .X(_07465_));
 sky130_fd_sc_hd__buf_4 _14852_ (.A(_07356_),
    .X(_07466_));
 sky130_fd_sc_hd__a22o_2 _14853_ (.A1(_07460_),
    .A2(_07461_),
    .B1(_07465_),
    .B2(_07466_),
    .X(_07467_));
 sky130_fd_sc_hd__clkbuf_4 _14854_ (.A(_07467_),
    .X(_07468_));
 sky130_fd_sc_hd__buf_2 _14855_ (.A(_07355_),
    .X(_07469_));
 sky130_fd_sc_hd__clkbuf_4 _14856_ (.A(_07435_),
    .X(_07470_));
 sky130_fd_sc_hd__buf_2 _14857_ (.A(_07443_),
    .X(_07471_));
 sky130_fd_sc_hd__clkbuf_4 _14858_ (.A(_07455_),
    .X(_07472_));
 sky130_fd_sc_hd__o22ai_1 _14859_ (.A1(_07470_),
    .A2(_07442_),
    .B1(_07471_),
    .B2(_07472_),
    .Y(_07473_));
 sky130_fd_sc_hd__or4bb_1 _14860_ (.A(_07468_),
    .B(_07469_),
    .C_N(_07456_),
    .D_N(_07473_),
    .X(_07474_));
 sky130_fd_sc_hd__nand2_1 _14861_ (.A(_07456_),
    .B(_07474_),
    .Y(_07475_));
 sky130_fd_sc_hd__or2b_1 _14862_ (.A(_07426_),
    .B_N(_07475_),
    .X(_07476_));
 sky130_fd_sc_hd__o22ai_1 _14863_ (.A1(_07378_),
    .A2(_07387_),
    .B1(_07399_),
    .B2(_07424_),
    .Y(_07477_));
 sky130_fd_sc_hd__a21o_1 _14864_ (.A1(_07100_),
    .A2(_07171_),
    .B1(_07336_),
    .X(_07478_));
 sky130_fd_sc_hd__mux2_1 _14865_ (.A0(_05093_),
    .A1(_05242_),
    .S(\rbzero.wall_tracer.side ),
    .X(_07479_));
 sky130_fd_sc_hd__nand2_1 _14866_ (.A(_07346_),
    .B(_07479_),
    .Y(_07480_));
 sky130_fd_sc_hd__a21o_2 _14867_ (.A1(_07478_),
    .A2(_07480_),
    .B1(_07349_),
    .X(_07481_));
 sky130_fd_sc_hd__a21oi_2 _14868_ (.A1(_07349_),
    .A2(\rbzero.wall_tracer.stepDistY[-7] ),
    .B1(\rbzero.wall_tracer.state[6] ),
    .Y(_07482_));
 sky130_fd_sc_hd__nor2_2 _14869_ (.A(_04927_),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .Y(_07483_));
 sky130_fd_sc_hd__a21o_1 _14870_ (.A1(_07481_),
    .A2(_07482_),
    .B1(_07483_),
    .X(_07484_));
 sky130_fd_sc_hd__buf_2 _14871_ (.A(_07484_),
    .X(_07485_));
 sky130_fd_sc_hd__nor2_1 _14872_ (.A(_07416_),
    .B(_07485_),
    .Y(_07486_));
 sky130_fd_sc_hd__or4_1 _14873_ (.A(_07378_),
    .B(_07387_),
    .C(_07399_),
    .D(_07423_),
    .X(_07487_));
 sky130_fd_sc_hd__a21bo_1 _14874_ (.A1(_07477_),
    .A2(_07486_),
    .B1_N(_07487_),
    .X(_07488_));
 sky130_fd_sc_hd__xnor2_1 _14875_ (.A(_07475_),
    .B(_07426_),
    .Y(_07489_));
 sky130_fd_sc_hd__nand2_1 _14876_ (.A(_07488_),
    .B(_07489_),
    .Y(_07490_));
 sky130_fd_sc_hd__buf_4 _14877_ (.A(_07374_),
    .X(_07491_));
 sky130_fd_sc_hd__or2_1 _14878_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_07411_),
    .X(_07492_));
 sky130_fd_sc_hd__inv_2 _14879_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .Y(_07493_));
 sky130_fd_sc_hd__inv_2 _14880_ (.A(\rbzero.debug_overlay.playerX[-1] ),
    .Y(_07494_));
 sky130_fd_sc_hd__and3b_1 _14881_ (.A_N(_07492_),
    .B(_07493_),
    .C(_07494_),
    .X(_07495_));
 sky130_fd_sc_hd__nand2_1 _14882_ (.A(\rbzero.wall_tracer.visualWallDist[0] ),
    .B(_03794_),
    .Y(_07496_));
 sky130_fd_sc_hd__or2_1 _14883_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .B(_07404_),
    .X(_07497_));
 sky130_fd_sc_hd__or3_1 _14884_ (.A(\rbzero.debug_overlay.playerY[-1] ),
    .B(\rbzero.debug_overlay.playerY[-2] ),
    .C(_07497_),
    .X(_07498_));
 sky130_fd_sc_hd__or3_1 _14885_ (.A(_03794_),
    .B(_05114_),
    .C(_07498_),
    .X(_07499_));
 sky130_fd_sc_hd__a21oi_2 _14886_ (.A1(_07496_),
    .A2(_07499_),
    .B1(_07466_),
    .Y(_07500_));
 sky130_fd_sc_hd__a31oi_4 _14887_ (.A1(_04937_),
    .A2(_07491_),
    .A3(_07495_),
    .B1(_07500_),
    .Y(_07501_));
 sky130_fd_sc_hd__a21o_1 _14888_ (.A1(_07213_),
    .A2(_07156_),
    .B1(_07346_),
    .X(_07502_));
 sky130_fd_sc_hd__o21a_1 _14889_ (.A1(_07341_),
    .A2(_05096_),
    .B1(_07336_),
    .X(_07503_));
 sky130_fd_sc_hd__o21ai_1 _14890_ (.A1(_07334_),
    .A2(_05258_),
    .B1(_07503_),
    .Y(_07504_));
 sky130_fd_sc_hd__a21o_1 _14891_ (.A1(_07502_),
    .A2(_07504_),
    .B1(_07351_),
    .X(_07505_));
 sky130_fd_sc_hd__a21oi_1 _14892_ (.A1(_07408_),
    .A2(\rbzero.wall_tracer.stepDistY[-9] ),
    .B1(_07352_),
    .Y(_07506_));
 sky130_fd_sc_hd__a2bb2o_2 _14893_ (.A1_N(_04928_),
    .A2_N(\rbzero.wall_tracer.stepDistX[-9] ),
    .B1(_07505_),
    .B2(_07506_),
    .X(_07507_));
 sky130_fd_sc_hd__buf_2 _14894_ (.A(_07507_),
    .X(_07508_));
 sky130_fd_sc_hd__nand2_4 _14895_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_03795_),
    .Y(_07509_));
 sky130_fd_sc_hd__or2_1 _14896_ (.A(_07466_),
    .B(_07509_),
    .X(_07510_));
 sky130_fd_sc_hd__nand2_1 _14897_ (.A(\rbzero.wall_tracer.state[13] ),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .Y(_07511_));
 sky130_fd_sc_hd__inv_2 _14898_ (.A(_07511_),
    .Y(_07512_));
 sky130_fd_sc_hd__mux2_1 _14899_ (.A0(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-2] ),
    .S(\rbzero.wall_tracer.side ),
    .X(_07513_));
 sky130_fd_sc_hd__o21ai_1 _14900_ (.A1(_04932_),
    .A2(_07513_),
    .B1(_03793_),
    .Y(_07514_));
 sky130_fd_sc_hd__a31o_2 _14901_ (.A1(_04932_),
    .A2(_07100_),
    .A3(_07146_),
    .B1(_07514_),
    .X(_07515_));
 sky130_fd_sc_hd__nand2_2 _14902_ (.A(_04928_),
    .B(_07515_),
    .Y(_07516_));
 sky130_fd_sc_hd__nor2_4 _14903_ (.A(_07512_),
    .B(_07516_),
    .Y(_07517_));
 sky130_fd_sc_hd__or4_1 _14904_ (.A(_07501_),
    .B(_07508_),
    .C(_07510_),
    .D(_07517_),
    .X(_07518_));
 sky130_fd_sc_hd__buf_4 _14905_ (.A(_04937_),
    .X(_07519_));
 sky130_fd_sc_hd__nor2_4 _14906_ (.A(_07519_),
    .B(_07509_),
    .Y(_07520_));
 sky130_fd_sc_hd__or3b_4 _14907_ (.A(_07352_),
    .B(_07512_),
    .C_N(_07515_),
    .X(_07521_));
 sky130_fd_sc_hd__a2bb2o_1 _14908_ (.A1_N(_07501_),
    .A2_N(_07508_),
    .B1(_07520_),
    .B2(_07521_),
    .X(_07522_));
 sky130_fd_sc_hd__nand2_1 _14909_ (.A(_07518_),
    .B(_07522_),
    .Y(_07523_));
 sky130_fd_sc_hd__nand2_2 _14910_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_03796_),
    .Y(_07524_));
 sky130_fd_sc_hd__inv_2 _14911_ (.A(\rbzero.wall_tracer.stepDistY[-11] ),
    .Y(_07525_));
 sky130_fd_sc_hd__a21o_1 _14912_ (.A1(_07100_),
    .A2(_07135_),
    .B1(_07336_),
    .X(_07526_));
 sky130_fd_sc_hd__mux2_1 _14913_ (.A0(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-3] ),
    .S(\rbzero.wall_tracer.side ),
    .X(_07527_));
 sky130_fd_sc_hd__a21oi_2 _14914_ (.A1(_07336_),
    .A2(_07527_),
    .B1(\rbzero.wall_tracer.state[13] ),
    .Y(_07528_));
 sky130_fd_sc_hd__a221o_4 _14915_ (.A1(_07349_),
    .A2(_07525_),
    .B1(_07526_),
    .B2(_07528_),
    .C1(_07352_),
    .X(_07529_));
 sky130_fd_sc_hd__or3_1 _14916_ (.A(_07523_),
    .B(_07524_),
    .C(_07529_),
    .X(_07530_));
 sky130_fd_sc_hd__o21ai_1 _14917_ (.A1(_07524_),
    .A2(_07529_),
    .B1(_07523_),
    .Y(_07531_));
 sky130_fd_sc_hd__and2_1 _14918_ (.A(_07530_),
    .B(_07531_),
    .X(_07532_));
 sky130_fd_sc_hd__nand2_1 _14919_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .B(_07404_),
    .Y(_07533_));
 sky130_fd_sc_hd__and2_1 _14920_ (.A(_07497_),
    .B(_07533_),
    .X(_07534_));
 sky130_fd_sc_hd__mux2_1 _14921_ (.A0(_07534_),
    .A1(\rbzero.debug_overlay.playerY[-3] ),
    .S(_05113_),
    .X(_07535_));
 sky130_fd_sc_hd__mux2_1 _14922_ (.A0(\rbzero.wall_tracer.visualWallDist[-3] ),
    .A1(_07535_),
    .S(_07349_),
    .X(_07536_));
 sky130_fd_sc_hd__inv_2 _14923_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .Y(_07537_));
 sky130_fd_sc_hd__nand2_1 _14924_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_07411_),
    .Y(_07538_));
 sky130_fd_sc_hd__nand2_1 _14925_ (.A(_07492_),
    .B(_07538_),
    .Y(_07539_));
 sky130_fd_sc_hd__mux2_1 _14926_ (.A0(_07537_),
    .A1(_07539_),
    .S(_07374_),
    .X(_07540_));
 sky130_fd_sc_hd__nand2_1 _14927_ (.A(_07356_),
    .B(_07540_),
    .Y(_07541_));
 sky130_fd_sc_hd__o21ai_4 _14928_ (.A1(_07356_),
    .A2(_07536_),
    .B1(_07541_),
    .Y(_07542_));
 sky130_fd_sc_hd__xor2_1 _14929_ (.A(\rbzero.debug_overlay.playerY[-2] ),
    .B(_07497_),
    .X(_07543_));
 sky130_fd_sc_hd__mux2_1 _14930_ (.A0(_07543_),
    .A1(\rbzero.debug_overlay.playerY[-2] ),
    .S(_05113_),
    .X(_07544_));
 sky130_fd_sc_hd__mux2_1 _14931_ (.A0(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A1(_07544_),
    .S(_07408_),
    .X(_07545_));
 sky130_fd_sc_hd__xnor2_1 _14932_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .B(_07492_),
    .Y(_07546_));
 sky130_fd_sc_hd__mux2_1 _14933_ (.A0(_07493_),
    .A1(_07546_),
    .S(_07374_),
    .X(_07547_));
 sky130_fd_sc_hd__nand2_1 _14934_ (.A(_07356_),
    .B(_07547_),
    .Y(_07548_));
 sky130_fd_sc_hd__o21ai_2 _14935_ (.A1(_04936_),
    .A2(_07545_),
    .B1(_07548_),
    .Y(_07549_));
 sky130_fd_sc_hd__clkbuf_4 _14936_ (.A(_07549_),
    .X(_07550_));
 sky130_fd_sc_hd__or4_1 _14937_ (.A(_07423_),
    .B(_07485_),
    .C(_07542_),
    .D(_07550_),
    .X(_07551_));
 sky130_fd_sc_hd__buf_2 _14938_ (.A(_07542_),
    .X(_07552_));
 sky130_fd_sc_hd__clkinv_4 _14939_ (.A(_07550_),
    .Y(_07553_));
 sky130_fd_sc_hd__a21oi_4 _14940_ (.A1(_07481_),
    .A2(_07482_),
    .B1(_07483_),
    .Y(_07554_));
 sky130_fd_sc_hd__a2bb2o_1 _14941_ (.A1_N(_07424_),
    .A2_N(_07552_),
    .B1(_07553_),
    .B2(_07554_),
    .X(_07555_));
 sky130_fd_sc_hd__nand2_1 _14942_ (.A(_07551_),
    .B(_07555_),
    .Y(_07556_));
 sky130_fd_sc_hd__o21ai_1 _14943_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_07497_),
    .B1(\rbzero.debug_overlay.playerY[-1] ),
    .Y(_07557_));
 sky130_fd_sc_hd__and2_1 _14944_ (.A(_07498_),
    .B(_07557_),
    .X(_07558_));
 sky130_fd_sc_hd__mux2_1 _14945_ (.A0(_07558_),
    .A1(\rbzero.debug_overlay.playerY[-1] ),
    .S(_05114_),
    .X(_07559_));
 sky130_fd_sc_hd__nand2_1 _14946_ (.A(_07453_),
    .B(_07559_),
    .Y(_07560_));
 sky130_fd_sc_hd__a21oi_1 _14947_ (.A1(\rbzero.wall_tracer.visualWallDist[-1] ),
    .A2(_03795_),
    .B1(_07466_),
    .Y(_07561_));
 sky130_fd_sc_hd__or3_1 _14948_ (.A(\rbzero.debug_overlay.playerX[-1] ),
    .B(\rbzero.debug_overlay.playerX[-2] ),
    .C(_07492_),
    .X(_07562_));
 sky130_fd_sc_hd__o21ai_1 _14949_ (.A1(\rbzero.debug_overlay.playerX[-2] ),
    .A2(_07492_),
    .B1(\rbzero.debug_overlay.playerX[-1] ),
    .Y(_07563_));
 sky130_fd_sc_hd__nand2_1 _14950_ (.A(_07562_),
    .B(_07563_),
    .Y(_07564_));
 sky130_fd_sc_hd__mux2_1 _14951_ (.A0(_07494_),
    .A1(_07564_),
    .S(_07374_),
    .X(_07565_));
 sky130_fd_sc_hd__a22o_1 _14952_ (.A1(_07560_),
    .A2(_07561_),
    .B1(_07565_),
    .B2(_04937_),
    .X(_07566_));
 sky130_fd_sc_hd__buf_2 _14953_ (.A(_07566_),
    .X(_07567_));
 sky130_fd_sc_hd__a21o_1 _14954_ (.A1(_07213_),
    .A2(_07164_),
    .B1(_07346_),
    .X(_07568_));
 sky130_fd_sc_hd__o21a_1 _14955_ (.A1(_07341_),
    .A2(_05095_),
    .B1(_07336_),
    .X(_07569_));
 sky130_fd_sc_hd__o21ai_1 _14956_ (.A1(_07334_),
    .A2(_05247_),
    .B1(_07569_),
    .Y(_07570_));
 sky130_fd_sc_hd__a21o_2 _14957_ (.A1(_07568_),
    .A2(_07570_),
    .B1(_07408_),
    .X(_07571_));
 sky130_fd_sc_hd__a21oi_4 _14958_ (.A1(_07408_),
    .A2(\rbzero.wall_tracer.stepDistY[-8] ),
    .B1(_07352_),
    .Y(_07572_));
 sky130_fd_sc_hd__nor2_2 _14959_ (.A(_04927_),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .Y(_07573_));
 sky130_fd_sc_hd__a21o_1 _14960_ (.A1(_07571_),
    .A2(_07572_),
    .B1(_07573_),
    .X(_07574_));
 sky130_fd_sc_hd__buf_2 _14961_ (.A(_07574_),
    .X(_07575_));
 sky130_fd_sc_hd__or2_1 _14962_ (.A(_07567_),
    .B(_07575_),
    .X(_07576_));
 sky130_fd_sc_hd__xnor2_1 _14963_ (.A(_07556_),
    .B(_07576_),
    .Y(_07577_));
 sky130_fd_sc_hd__or4_1 _14964_ (.A(_07485_),
    .B(_07542_),
    .C(_07550_),
    .D(_07575_),
    .X(_07578_));
 sky130_fd_sc_hd__a21oi_4 _14965_ (.A1(_07571_),
    .A2(_07572_),
    .B1(_07573_),
    .Y(_07579_));
 sky130_fd_sc_hd__a2bb2o_1 _14966_ (.A1_N(_07485_),
    .A2_N(_07552_),
    .B1(_07553_),
    .B2(_07579_),
    .X(_07580_));
 sky130_fd_sc_hd__nand2_1 _14967_ (.A(_07578_),
    .B(_07580_),
    .Y(_07581_));
 sky130_fd_sc_hd__or2_1 _14968_ (.A(_07508_),
    .B(_07567_),
    .X(_07582_));
 sky130_fd_sc_hd__o21a_1 _14969_ (.A1(_07581_),
    .A2(_07582_),
    .B1(_07578_),
    .X(_07583_));
 sky130_fd_sc_hd__nor2_1 _14970_ (.A(_07577_),
    .B(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__nand2_1 _14971_ (.A(_07577_),
    .B(_07583_),
    .Y(_07585_));
 sky130_fd_sc_hd__and2b_1 _14972_ (.A_N(_07584_),
    .B(_07585_),
    .X(_07586_));
 sky130_fd_sc_hd__xnor2_1 _14973_ (.A(_07532_),
    .B(_07586_),
    .Y(_07587_));
 sky130_fd_sc_hd__a21o_1 _14974_ (.A1(_07476_),
    .A2(_07490_),
    .B1(_07587_),
    .X(_07588_));
 sky130_fd_sc_hd__nand3_1 _14975_ (.A(_07476_),
    .B(_07490_),
    .C(_07587_),
    .Y(_07589_));
 sky130_fd_sc_hd__nand2_1 _14976_ (.A(_07588_),
    .B(_07589_),
    .Y(_07590_));
 sky130_fd_sc_hd__buf_2 _14977_ (.A(_07501_),
    .X(_07591_));
 sky130_fd_sc_hd__o21ai_4 _14978_ (.A1(_04928_),
    .A2(\rbzero.wall_tracer.stepDistX[-10] ),
    .B1(_07521_),
    .Y(_07592_));
 sky130_fd_sc_hd__buf_2 _14979_ (.A(_07592_),
    .X(_07593_));
 sky130_fd_sc_hd__nor2_1 _14980_ (.A(_07591_),
    .B(_07593_),
    .Y(_07594_));
 sky130_fd_sc_hd__nor2_1 _14981_ (.A(_07509_),
    .B(_07529_),
    .Y(_07595_));
 sky130_fd_sc_hd__xnor2_1 _14982_ (.A(_07594_),
    .B(_07595_),
    .Y(_07596_));
 sky130_fd_sc_hd__or2_1 _14983_ (.A(_07519_),
    .B(_07524_),
    .X(_07597_));
 sky130_fd_sc_hd__buf_2 _14984_ (.A(_07597_),
    .X(_07598_));
 sky130_fd_sc_hd__a21o_1 _14985_ (.A1(_07213_),
    .A2(_07117_),
    .B1(_07346_),
    .X(_07599_));
 sky130_fd_sc_hd__mux2_1 _14986_ (.A0(\rbzero.wall_tracer.rayAddendY[-4] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-4] ),
    .S(_07341_),
    .X(_07600_));
 sky130_fd_sc_hd__a21oi_2 _14987_ (.A1(_07346_),
    .A2(_07600_),
    .B1(_07349_),
    .Y(_07601_));
 sky130_fd_sc_hd__and2_2 _14988_ (.A(_07599_),
    .B(_07601_),
    .X(_07602_));
 sky130_fd_sc_hd__nor2_1 _14989_ (.A(_07598_),
    .B(_07602_),
    .Y(_07603_));
 sky130_fd_sc_hd__xnor2_1 _14990_ (.A(_07596_),
    .B(_07603_),
    .Y(_07604_));
 sky130_fd_sc_hd__xnor2_1 _14991_ (.A(_07581_),
    .B(_07582_),
    .Y(_07605_));
 sky130_fd_sc_hd__or4_1 _14992_ (.A(_07507_),
    .B(_07542_),
    .C(_07549_),
    .D(_07575_),
    .X(_07606_));
 sky130_fd_sc_hd__inv_2 _14993_ (.A(_07606_),
    .Y(_07607_));
 sky130_fd_sc_hd__o22ai_1 _14994_ (.A1(_07508_),
    .A2(_07550_),
    .B1(_07575_),
    .B2(_07542_),
    .Y(_07608_));
 sky130_fd_sc_hd__nor2_1 _14995_ (.A(_07566_),
    .B(_07593_),
    .Y(_07609_));
 sky130_fd_sc_hd__and3_1 _14996_ (.A(_07606_),
    .B(_07608_),
    .C(_07609_),
    .X(_07610_));
 sky130_fd_sc_hd__nor2_1 _14997_ (.A(_07607_),
    .B(_07610_),
    .Y(_07611_));
 sky130_fd_sc_hd__nand2_1 _14998_ (.A(_07605_),
    .B(_07611_),
    .Y(_07612_));
 sky130_fd_sc_hd__nor2_1 _14999_ (.A(_07605_),
    .B(_07611_),
    .Y(_07613_));
 sky130_fd_sc_hd__a21o_1 _15000_ (.A1(_07604_),
    .A2(_07612_),
    .B1(_07613_),
    .X(_07614_));
 sky130_fd_sc_hd__or2b_1 _15001_ (.A(_07590_),
    .B_N(_07614_),
    .X(_07615_));
 sky130_fd_sc_hd__a21o_4 _15002_ (.A1(_07526_),
    .A2(_07528_),
    .B1(_07356_),
    .X(_07616_));
 sky130_fd_sc_hd__nand2_1 _15003_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_03796_),
    .Y(_07617_));
 sky130_fd_sc_hd__buf_2 _15004_ (.A(_07617_),
    .X(_07618_));
 sky130_fd_sc_hd__nand2_4 _15005_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_03796_),
    .Y(_07619_));
 sky130_fd_sc_hd__or2_2 _15006_ (.A(_07519_),
    .B(_07619_),
    .X(_07620_));
 sky130_fd_sc_hd__buf_2 _15007_ (.A(_07620_),
    .X(_07621_));
 sky130_fd_sc_hd__or2_1 _15008_ (.A(_07602_),
    .B(_07621_),
    .X(_07622_));
 sky130_fd_sc_hd__nor3_1 _15009_ (.A(_07616_),
    .B(_07618_),
    .C(_07622_),
    .Y(_07623_));
 sky130_fd_sc_hd__or2_1 _15010_ (.A(_07519_),
    .B(_07602_),
    .X(_07624_));
 sky130_fd_sc_hd__buf_2 _15011_ (.A(_07624_),
    .X(_07625_));
 sky130_fd_sc_hd__o22a_1 _15012_ (.A1(_07616_),
    .A2(_07619_),
    .B1(_07618_),
    .B2(_07625_),
    .X(_07626_));
 sky130_fd_sc_hd__or2_1 _15013_ (.A(_07623_),
    .B(_07626_),
    .X(_07627_));
 sky130_fd_sc_hd__a21o_1 _15014_ (.A1(_07518_),
    .A2(_07530_),
    .B1(_07627_),
    .X(_07628_));
 sky130_fd_sc_hd__nand3_1 _15015_ (.A(_07518_),
    .B(_07530_),
    .C(_07627_),
    .Y(_07629_));
 sky130_fd_sc_hd__and2_1 _15016_ (.A(_07628_),
    .B(_07629_),
    .X(_07630_));
 sky130_fd_sc_hd__clkbuf_4 _15017_ (.A(_07524_),
    .X(_07631_));
 sky130_fd_sc_hd__a21oi_4 _15018_ (.A1(_07599_),
    .A2(_07601_),
    .B1(_07352_),
    .Y(_07632_));
 sky130_fd_sc_hd__o21ai_4 _15019_ (.A1(_03794_),
    .A2(\rbzero.wall_tracer.stepDistY[-12] ),
    .B1(_07632_),
    .Y(_07633_));
 sky130_fd_sc_hd__nand2_1 _15020_ (.A(_07594_),
    .B(_07595_),
    .Y(_07634_));
 sky130_fd_sc_hd__o31a_1 _15021_ (.A1(_07631_),
    .A2(_07596_),
    .A3(_07633_),
    .B1(_07634_),
    .X(_07635_));
 sky130_fd_sc_hd__nor2_1 _15022_ (.A(_07622_),
    .B(_07635_),
    .Y(_07636_));
 sky130_fd_sc_hd__nand2_1 _15023_ (.A(_07630_),
    .B(_07636_),
    .Y(_07637_));
 sky130_fd_sc_hd__or2_1 _15024_ (.A(_07630_),
    .B(_07636_),
    .X(_07638_));
 sky130_fd_sc_hd__nand2_1 _15025_ (.A(_07637_),
    .B(_07638_),
    .Y(_07639_));
 sky130_fd_sc_hd__a21oi_2 _15026_ (.A1(_07588_),
    .A2(_07615_),
    .B1(_07639_),
    .Y(_07640_));
 sky130_fd_sc_hd__nand2_1 _15027_ (.A(_07466_),
    .B(\rbzero.wall_tracer.stepDistX[1] ),
    .Y(_07641_));
 sky130_fd_sc_hd__or2_1 _15028_ (.A(\rbzero.wall_tracer.visualWallDist[-9] ),
    .B(\rbzero.wall_tracer.state[13] ),
    .X(_07642_));
 sky130_fd_sc_hd__o211a_1 _15029_ (.A1(\rbzero.debug_overlay.playerY[-9] ),
    .A2(_03793_),
    .B1(_04927_),
    .C1(_07642_),
    .X(_07643_));
 sky130_fd_sc_hd__a21oi_1 _15030_ (.A1(\rbzero.debug_overlay.playerX[-9] ),
    .A2(\rbzero.wall_tracer.state[6] ),
    .B1(_07643_),
    .Y(_07644_));
 sky130_fd_sc_hd__clkbuf_4 _15031_ (.A(_07644_),
    .X(_07645_));
 sky130_fd_sc_hd__clkbuf_4 _15032_ (.A(_07645_),
    .X(_07646_));
 sky130_fd_sc_hd__a21oi_1 _15033_ (.A1(_07455_),
    .A2(_07641_),
    .B1(_07646_),
    .Y(_07647_));
 sky130_fd_sc_hd__xnor2_4 _15034_ (.A(_07208_),
    .B(_07445_),
    .Y(_07648_));
 sky130_fd_sc_hd__mux2_1 _15035_ (.A0(_05106_),
    .A1(_05273_),
    .S(_07342_),
    .X(_07649_));
 sky130_fd_sc_hd__a21o_1 _15036_ (.A1(_07337_),
    .A2(_07649_),
    .B1(_07408_),
    .X(_07650_));
 sky130_fd_sc_hd__a21o_4 _15037_ (.A1(_04933_),
    .A2(_07648_),
    .B1(_07650_),
    .X(_07651_));
 sky130_fd_sc_hd__nor2_2 _15038_ (.A(_07260_),
    .B(_07351_),
    .Y(_07652_));
 sky130_fd_sc_hd__and3_1 _15039_ (.A(_04928_),
    .B(_07651_),
    .C(_07652_),
    .X(_07653_));
 sky130_fd_sc_hd__xnor2_1 _15040_ (.A(_07647_),
    .B(_07653_),
    .Y(_07654_));
 sky130_fd_sc_hd__and2_1 _15041_ (.A(_07100_),
    .B(_07210_),
    .X(_07655_));
 sky130_fd_sc_hd__a31o_1 _15042_ (.A1(_07028_),
    .A2(_07076_),
    .A3(_07098_),
    .B1(_07133_),
    .X(_07656_));
 sky130_fd_sc_hd__o211a_1 _15043_ (.A1(_07446_),
    .A2(_07448_),
    .B1(_07656_),
    .C1(_07447_),
    .X(_07657_));
 sky130_fd_sc_hd__xnor2_2 _15044_ (.A(_07655_),
    .B(_07657_),
    .Y(_07658_));
 sky130_fd_sc_hd__nand2_1 _15045_ (.A(_07342_),
    .B(_05196_),
    .Y(_07659_));
 sky130_fd_sc_hd__o211a_1 _15046_ (.A1(_07342_),
    .A2(_05073_),
    .B1(_07659_),
    .C1(_07337_),
    .X(_07660_));
 sky130_fd_sc_hd__a211o_1 _15047_ (.A1(_04932_),
    .A2(_07658_),
    .B1(_07660_),
    .C1(_07453_),
    .X(_07661_));
 sky130_fd_sc_hd__o21a_1 _15048_ (.A1(_03795_),
    .A2(\rbzero.wall_tracer.stepDistY[3] ),
    .B1(_04928_),
    .X(_07662_));
 sky130_fd_sc_hd__nand2_4 _15049_ (.A(_07661_),
    .B(_07662_),
    .Y(_07663_));
 sky130_fd_sc_hd__nand2_4 _15050_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_03793_),
    .Y(_07664_));
 sky130_fd_sc_hd__nor2_1 _15051_ (.A(_07663_),
    .B(_07664_),
    .Y(_07665_));
 sky130_fd_sc_hd__xor2_1 _15052_ (.A(_07654_),
    .B(_07665_),
    .X(_07666_));
 sky130_fd_sc_hd__xnor2_2 _15053_ (.A(_07202_),
    .B(_07448_),
    .Y(_07667_));
 sky130_fd_sc_hd__nor2_1 _15054_ (.A(_07341_),
    .B(_05110_),
    .Y(_07668_));
 sky130_fd_sc_hd__a211o_1 _15055_ (.A1(_07342_),
    .A2(_05267_),
    .B1(_07668_),
    .C1(_04932_),
    .X(_07669_));
 sky130_fd_sc_hd__o21ai_4 _15056_ (.A1(_07337_),
    .A2(_07667_),
    .B1(_07669_),
    .Y(_07670_));
 sky130_fd_sc_hd__nor2_1 _15057_ (.A(_03794_),
    .B(\rbzero.wall_tracer.stepDistY[0] ),
    .Y(_07671_));
 sky130_fd_sc_hd__a211o_2 _15058_ (.A1(_03794_),
    .A2(_07670_),
    .B1(_07671_),
    .C1(_07356_),
    .X(_07672_));
 sky130_fd_sc_hd__nand2_2 _15059_ (.A(_04936_),
    .B(\rbzero.wall_tracer.stepDistX[0] ),
    .Y(_07673_));
 sky130_fd_sc_hd__a21o_1 _15060_ (.A1(_07672_),
    .A2(_07673_),
    .B1(_07646_),
    .X(_07674_));
 sky130_fd_sc_hd__nand2_2 _15061_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_03794_),
    .Y(_07675_));
 sky130_fd_sc_hd__nor2_1 _15062_ (.A(_07455_),
    .B(_07675_),
    .Y(_07676_));
 sky130_fd_sc_hd__xnor2_1 _15063_ (.A(_07674_),
    .B(_07676_),
    .Y(_07677_));
 sky130_fd_sc_hd__nand2_1 _15064_ (.A(_04929_),
    .B(_07651_),
    .Y(_07678_));
 sky130_fd_sc_hd__nor2_1 _15065_ (.A(_07678_),
    .B(_07664_),
    .Y(_07679_));
 sky130_fd_sc_hd__clkbuf_4 _15066_ (.A(_07675_),
    .X(_07680_));
 sky130_fd_sc_hd__or3_1 _15067_ (.A(_07472_),
    .B(_07680_),
    .C(_07674_),
    .X(_07681_));
 sky130_fd_sc_hd__a21boi_1 _15068_ (.A1(_07677_),
    .A2(_07679_),
    .B1_N(_07681_),
    .Y(_07682_));
 sky130_fd_sc_hd__xor2_1 _15069_ (.A(_07666_),
    .B(_07682_),
    .X(_07683_));
 sky130_fd_sc_hd__and2_1 _15070_ (.A(_07672_),
    .B(_07673_),
    .X(_07684_));
 sky130_fd_sc_hd__buf_2 _15071_ (.A(_07684_),
    .X(_07685_));
 sky130_fd_sc_hd__and2_1 _15072_ (.A(_07453_),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .X(_07686_));
 sky130_fd_sc_hd__a2111o_1 _15073_ (.A1(_07202_),
    .A2(_07444_),
    .B1(_07211_),
    .C1(_07208_),
    .D1(_07206_),
    .X(_07687_));
 sky130_fd_sc_hd__nor2_1 _15074_ (.A(_07217_),
    .B(_07687_),
    .Y(_07688_));
 sky130_fd_sc_hd__and2_1 _15075_ (.A(_07101_),
    .B(_07216_),
    .X(_07689_));
 sky130_fd_sc_hd__o2111a_1 _15076_ (.A1(_07446_),
    .A2(_07448_),
    .B1(_07655_),
    .C1(_07656_),
    .D1(_07447_),
    .X(_07690_));
 sky130_fd_sc_hd__nor2_1 _15077_ (.A(_07689_),
    .B(_07690_),
    .Y(_07691_));
 sky130_fd_sc_hd__a31o_1 _15078_ (.A1(_07334_),
    .A2(_05069_),
    .A3(_05112_),
    .B1(_04932_),
    .X(_07692_));
 sky130_fd_sc_hd__a21o_1 _15079_ (.A1(_07342_),
    .A2(_05186_),
    .B1(_07692_),
    .X(_07693_));
 sky130_fd_sc_hd__and2_4 _15080_ (.A(_03794_),
    .B(_07693_),
    .X(_07694_));
 sky130_fd_sc_hd__o31a_2 _15081_ (.A1(_07337_),
    .A2(_07688_),
    .A3(_07691_),
    .B1(_07694_),
    .X(_07695_));
 sky130_fd_sc_hd__o21ai_4 _15082_ (.A1(_07686_),
    .A2(_07695_),
    .B1(_04928_),
    .Y(_07696_));
 sky130_fd_sc_hd__clkinv_4 _15083_ (.A(_07434_),
    .Y(_07697_));
 sky130_fd_sc_hd__and2_4 _15084_ (.A(\rbzero.wall_tracer.visualWallDist[-12] ),
    .B(_03794_),
    .X(_07698_));
 sky130_fd_sc_hd__and4bb_1 _15085_ (.A_N(_07685_),
    .B_N(_07696_),
    .C(_07697_),
    .D(_07698_),
    .X(_07699_));
 sky130_fd_sc_hd__o22a_1 _15086_ (.A1(_07470_),
    .A2(_07685_),
    .B1(_07696_),
    .B2(_07471_),
    .X(_07700_));
 sky130_fd_sc_hd__or2_1 _15087_ (.A(_07699_),
    .B(_07700_),
    .X(_07701_));
 sky130_fd_sc_hd__inv_2 _15088_ (.A(\rbzero.wall_tracer.stepDistY[-1] ),
    .Y(_07702_));
 sky130_fd_sc_hd__o21a_1 _15089_ (.A1(_07195_),
    .A2(_07198_),
    .B1(_07213_),
    .X(_07703_));
 sky130_fd_sc_hd__a21o_1 _15090_ (.A1(_07444_),
    .A2(_07703_),
    .B1(_07337_),
    .X(_07704_));
 sky130_fd_sc_hd__nand2_1 _15091_ (.A(_07341_),
    .B(_05215_),
    .Y(_07705_));
 sky130_fd_sc_hd__o211a_1 _15092_ (.A1(_07342_),
    .A2(_05100_),
    .B1(_07705_),
    .C1(_07346_),
    .X(_07706_));
 sky130_fd_sc_hd__nor2_1 _15093_ (.A(_07351_),
    .B(_07706_),
    .Y(_07707_));
 sky130_fd_sc_hd__a221o_1 _15094_ (.A1(_07408_),
    .A2(_07702_),
    .B1(_07704_),
    .B2(_07707_),
    .C1(_04935_),
    .X(_07708_));
 sky130_fd_sc_hd__clkbuf_4 _15095_ (.A(_07708_),
    .X(_07709_));
 sky130_fd_sc_hd__nand2_1 _15096_ (.A(_07466_),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .Y(_07710_));
 sky130_fd_sc_hd__and2_1 _15097_ (.A(_07709_),
    .B(_07710_),
    .X(_07711_));
 sky130_fd_sc_hd__clkbuf_4 _15098_ (.A(_07711_),
    .X(_07712_));
 sky130_fd_sc_hd__nor2_1 _15099_ (.A(_07468_),
    .B(_07712_),
    .Y(_07713_));
 sky130_fd_sc_hd__xnor2_1 _15100_ (.A(_07701_),
    .B(_07713_),
    .Y(_07714_));
 sky130_fd_sc_hd__xnor2_1 _15101_ (.A(_07683_),
    .B(_07714_),
    .Y(_07715_));
 sky130_fd_sc_hd__xnor2_1 _15102_ (.A(_07677_),
    .B(_07679_),
    .Y(_07716_));
 sky130_fd_sc_hd__a21oi_1 _15103_ (.A1(_07709_),
    .A2(_07710_),
    .B1(_07646_),
    .Y(_07717_));
 sky130_fd_sc_hd__nand2_2 _15104_ (.A(_04927_),
    .B(_07652_),
    .Y(_07718_));
 sky130_fd_sc_hd__nor2_1 _15105_ (.A(_07670_),
    .B(_07718_),
    .Y(_07719_));
 sky130_fd_sc_hd__xor2_1 _15106_ (.A(_07717_),
    .B(_07719_),
    .X(_07720_));
 sky130_fd_sc_hd__nor2_1 _15107_ (.A(_07472_),
    .B(_07664_),
    .Y(_07721_));
 sky130_fd_sc_hd__nand2_1 _15108_ (.A(_07720_),
    .B(_07721_),
    .Y(_07722_));
 sky130_fd_sc_hd__a21boi_1 _15109_ (.A1(_07717_),
    .A2(_07719_),
    .B1_N(_07722_),
    .Y(_07723_));
 sky130_fd_sc_hd__xor2_1 _15110_ (.A(_07716_),
    .B(_07723_),
    .X(_07724_));
 sky130_fd_sc_hd__or4_1 _15111_ (.A(_07470_),
    .B(_07443_),
    .C(_07663_),
    .D(_07711_),
    .X(_07725_));
 sky130_fd_sc_hd__nand2_1 _15112_ (.A(_07709_),
    .B(_07710_),
    .Y(_07726_));
 sky130_fd_sc_hd__a32o_1 _15113_ (.A1(_07698_),
    .A2(_07661_),
    .A3(_07662_),
    .B1(_07726_),
    .B2(_07697_),
    .X(_07727_));
 sky130_fd_sc_hd__nand2_1 _15114_ (.A(_07725_),
    .B(_07727_),
    .Y(_07728_));
 sky130_fd_sc_hd__nor2_1 _15115_ (.A(_03794_),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .Y(_07729_));
 sky130_fd_sc_hd__a21o_1 _15116_ (.A1(_07213_),
    .A2(_07195_),
    .B1(_07346_),
    .X(_07730_));
 sky130_fd_sc_hd__nor2_1 _15117_ (.A(_07334_),
    .B(_05210_),
    .Y(_07731_));
 sky130_fd_sc_hd__a211o_1 _15118_ (.A1(_07334_),
    .A2(_05078_),
    .B1(_07731_),
    .C1(_04932_),
    .X(_07732_));
 sky130_fd_sc_hd__a21oi_1 _15119_ (.A1(_07730_),
    .A2(_07732_),
    .B1(_07351_),
    .Y(_07733_));
 sky130_fd_sc_hd__nand2_1 _15120_ (.A(_04935_),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .Y(_07734_));
 sky130_fd_sc_hd__o31a_2 _15121_ (.A1(_04935_),
    .A2(_07729_),
    .A3(_07733_),
    .B1(_07734_),
    .X(_07735_));
 sky130_fd_sc_hd__buf_2 _15122_ (.A(_07735_),
    .X(_07736_));
 sky130_fd_sc_hd__nor2_1 _15123_ (.A(_07468_),
    .B(_07736_),
    .Y(_07737_));
 sky130_fd_sc_hd__xnor2_1 _15124_ (.A(_07728_),
    .B(_07737_),
    .Y(_07738_));
 sky130_fd_sc_hd__nor2_1 _15125_ (.A(_07716_),
    .B(_07723_),
    .Y(_07739_));
 sky130_fd_sc_hd__a21oi_1 _15126_ (.A1(_07724_),
    .A2(_07738_),
    .B1(_07739_),
    .Y(_07740_));
 sky130_fd_sc_hd__xor2_1 _15127_ (.A(_07715_),
    .B(_07740_),
    .X(_07741_));
 sky130_fd_sc_hd__buf_2 _15128_ (.A(_07442_),
    .X(_07742_));
 sky130_fd_sc_hd__nor2_1 _15129_ (.A(_07742_),
    .B(_07400_),
    .Y(_07743_));
 sky130_fd_sc_hd__o22ai_1 _15130_ (.A1(_07442_),
    .A2(_07379_),
    .B1(_07400_),
    .B2(_07355_),
    .Y(_07744_));
 sky130_fd_sc_hd__nor2_1 _15131_ (.A(_07388_),
    .B(_07416_),
    .Y(_07745_));
 sky130_fd_sc_hd__a22oi_2 _15132_ (.A1(_07380_),
    .A2(_07743_),
    .B1(_07744_),
    .B2(_07745_),
    .Y(_07746_));
 sky130_fd_sc_hd__a21bo_1 _15133_ (.A1(_07727_),
    .A2(_07737_),
    .B1_N(_07725_),
    .X(_07747_));
 sky130_fd_sc_hd__nor2_1 _15134_ (.A(_07379_),
    .B(_07736_),
    .Y(_07748_));
 sky130_fd_sc_hd__or4_1 _15135_ (.A(_07442_),
    .B(_07379_),
    .C(_07399_),
    .D(_07735_),
    .X(_07749_));
 sky130_fd_sc_hd__o21ai_1 _15136_ (.A1(_07748_),
    .A2(_07743_),
    .B1(_07749_),
    .Y(_07750_));
 sky130_fd_sc_hd__clkbuf_4 _15137_ (.A(_07416_),
    .X(_07751_));
 sky130_fd_sc_hd__nor2_1 _15138_ (.A(_07469_),
    .B(_07751_),
    .Y(_07752_));
 sky130_fd_sc_hd__xnor2_1 _15139_ (.A(_07750_),
    .B(_07752_),
    .Y(_07753_));
 sky130_fd_sc_hd__xor2_1 _15140_ (.A(_07747_),
    .B(_07753_),
    .X(_07754_));
 sky130_fd_sc_hd__xnor2_1 _15141_ (.A(_07746_),
    .B(_07754_),
    .Y(_07755_));
 sky130_fd_sc_hd__xnor2_1 _15142_ (.A(_07741_),
    .B(_07755_),
    .Y(_07756_));
 sky130_fd_sc_hd__xnor2_1 _15143_ (.A(_07724_),
    .B(_07738_),
    .Y(_07757_));
 sky130_fd_sc_hd__xnor2_1 _15144_ (.A(_07720_),
    .B(_07721_),
    .Y(_07758_));
 sky130_fd_sc_hd__or4_1 _15145_ (.A(_07645_),
    .B(_07675_),
    .C(_07708_),
    .D(_07735_),
    .X(_07759_));
 sky130_fd_sc_hd__a21o_2 _15146_ (.A1(_03795_),
    .A2(_07670_),
    .B1(_07466_),
    .X(_07760_));
 sky130_fd_sc_hd__o22ai_1 _15147_ (.A1(_07675_),
    .A2(_07709_),
    .B1(_07735_),
    .B2(_07646_),
    .Y(_07761_));
 sky130_fd_sc_hd__or4bb_1 _15148_ (.A(_07760_),
    .B(_07664_),
    .C_N(_07759_),
    .D_N(_07761_),
    .X(_07762_));
 sky130_fd_sc_hd__and2_1 _15149_ (.A(_07759_),
    .B(_07762_),
    .X(_07763_));
 sky130_fd_sc_hd__xor2_1 _15150_ (.A(_07758_),
    .B(_07763_),
    .X(_07764_));
 sky130_fd_sc_hd__nor2_1 _15151_ (.A(_07470_),
    .B(_07735_),
    .Y(_07765_));
 sky130_fd_sc_hd__and4_1 _15152_ (.A(_04929_),
    .B(_07698_),
    .C(_07651_),
    .D(_07765_),
    .X(_07766_));
 sky130_fd_sc_hd__a31o_1 _15153_ (.A1(_04929_),
    .A2(_07698_),
    .A3(_07651_),
    .B1(_07765_),
    .X(_07767_));
 sky130_fd_sc_hd__and2b_1 _15154_ (.A_N(_07766_),
    .B(_07767_),
    .X(_07768_));
 sky130_fd_sc_hd__nor2_1 _15155_ (.A(_07742_),
    .B(_07468_),
    .Y(_07769_));
 sky130_fd_sc_hd__xor2_1 _15156_ (.A(_07768_),
    .B(_07769_),
    .X(_07770_));
 sky130_fd_sc_hd__nor2_1 _15157_ (.A(_07758_),
    .B(_07763_),
    .Y(_07771_));
 sky130_fd_sc_hd__a21oi_1 _15158_ (.A1(_07764_),
    .A2(_07770_),
    .B1(_07771_),
    .Y(_07772_));
 sky130_fd_sc_hd__xor2_1 _15159_ (.A(_07757_),
    .B(_07772_),
    .X(_07773_));
 sky130_fd_sc_hd__o31a_1 _15160_ (.A1(_07403_),
    .A2(_07751_),
    .A3(_07424_),
    .B1(_07402_),
    .X(_07774_));
 sky130_fd_sc_hd__a21o_1 _15161_ (.A1(_07767_),
    .A2(_07769_),
    .B1(_07766_),
    .X(_07775_));
 sky130_fd_sc_hd__a21boi_1 _15162_ (.A1(_07380_),
    .A2(_07743_),
    .B1_N(_07744_),
    .Y(_07776_));
 sky130_fd_sc_hd__xnor2_1 _15163_ (.A(_07776_),
    .B(_07745_),
    .Y(_07777_));
 sky130_fd_sc_hd__xnor2_1 _15164_ (.A(_07775_),
    .B(_07777_),
    .Y(_07778_));
 sky130_fd_sc_hd__xnor2_1 _15165_ (.A(_07774_),
    .B(_07778_),
    .Y(_07779_));
 sky130_fd_sc_hd__nor2_1 _15166_ (.A(_07757_),
    .B(_07772_),
    .Y(_07780_));
 sky130_fd_sc_hd__a21oi_1 _15167_ (.A1(_07773_),
    .A2(_07779_),
    .B1(_07780_),
    .Y(_07781_));
 sky130_fd_sc_hd__nor2_1 _15168_ (.A(_07756_),
    .B(_07781_),
    .Y(_07782_));
 sky130_fd_sc_hd__xor2_1 _15169_ (.A(_07756_),
    .B(_07781_),
    .X(_07783_));
 sky130_fd_sc_hd__a21o_1 _15170_ (.A1(_07532_),
    .A2(_07585_),
    .B1(_07584_),
    .X(_07784_));
 sky130_fd_sc_hd__or2b_1 _15171_ (.A(_07777_),
    .B_N(_07775_),
    .X(_07785_));
 sky130_fd_sc_hd__or2b_1 _15172_ (.A(_07774_),
    .B_N(_07778_),
    .X(_07786_));
 sky130_fd_sc_hd__nand2_1 _15173_ (.A(_07785_),
    .B(_07786_),
    .Y(_07787_));
 sky130_fd_sc_hd__clkbuf_4 _15174_ (.A(_07517_),
    .X(_07788_));
 sky130_fd_sc_hd__and2_1 _15175_ (.A(_07505_),
    .B(_07506_),
    .X(_07789_));
 sky130_fd_sc_hd__buf_2 _15176_ (.A(_07510_),
    .X(_07790_));
 sky130_fd_sc_hd__or4_1 _15177_ (.A(_07501_),
    .B(_07789_),
    .C(_07790_),
    .D(_07575_),
    .X(_07791_));
 sky130_fd_sc_hd__buf_2 _15178_ (.A(_07789_),
    .X(_07792_));
 sky130_fd_sc_hd__a31o_2 _15179_ (.A1(_07519_),
    .A2(_07491_),
    .A3(_07495_),
    .B1(_07500_),
    .X(_07793_));
 sky130_fd_sc_hd__a2bb2o_1 _15180_ (.A1_N(_07792_),
    .A2_N(_07790_),
    .B1(_07579_),
    .B2(_07793_),
    .X(_07794_));
 sky130_fd_sc_hd__nand2_1 _15181_ (.A(_07791_),
    .B(_07794_),
    .Y(_07795_));
 sky130_fd_sc_hd__or3_1 _15182_ (.A(_07788_),
    .B(_07598_),
    .C(_07795_),
    .X(_07796_));
 sky130_fd_sc_hd__o21ai_1 _15183_ (.A1(_07788_),
    .A2(_07598_),
    .B1(_07795_),
    .Y(_07797_));
 sky130_fd_sc_hd__and2_1 _15184_ (.A(_07796_),
    .B(_07797_),
    .X(_07798_));
 sky130_fd_sc_hd__or4_1 _15185_ (.A(_07387_),
    .B(_07424_),
    .C(_07552_),
    .D(_07550_),
    .X(_07799_));
 sky130_fd_sc_hd__buf_2 _15186_ (.A(_07550_),
    .X(_07800_));
 sky130_fd_sc_hd__o22ai_1 _15187_ (.A1(_07388_),
    .A2(_07552_),
    .B1(_07800_),
    .B2(_07424_),
    .Y(_07801_));
 sky130_fd_sc_hd__nand2_1 _15188_ (.A(_07799_),
    .B(_07801_),
    .Y(_07802_));
 sky130_fd_sc_hd__or2_1 _15189_ (.A(_07485_),
    .B(_07567_),
    .X(_07803_));
 sky130_fd_sc_hd__xnor2_1 _15190_ (.A(_07802_),
    .B(_07803_),
    .Y(_07804_));
 sky130_fd_sc_hd__clkbuf_4 _15191_ (.A(_07567_),
    .X(_07805_));
 sky130_fd_sc_hd__o31a_1 _15192_ (.A1(_07556_),
    .A2(_07805_),
    .A3(_07575_),
    .B1(_07551_),
    .X(_07806_));
 sky130_fd_sc_hd__nor2_1 _15193_ (.A(_07804_),
    .B(_07806_),
    .Y(_07807_));
 sky130_fd_sc_hd__nand2_1 _15194_ (.A(_07804_),
    .B(_07806_),
    .Y(_07808_));
 sky130_fd_sc_hd__and2b_1 _15195_ (.A_N(_07807_),
    .B(_07808_),
    .X(_07809_));
 sky130_fd_sc_hd__xnor2_1 _15196_ (.A(_07798_),
    .B(_07809_),
    .Y(_07810_));
 sky130_fd_sc_hd__xor2_1 _15197_ (.A(_07787_),
    .B(_07810_),
    .X(_07811_));
 sky130_fd_sc_hd__xnor2_1 _15198_ (.A(_07784_),
    .B(_07811_),
    .Y(_07812_));
 sky130_fd_sc_hd__and2_1 _15199_ (.A(_07783_),
    .B(_07812_),
    .X(_07813_));
 sky130_fd_sc_hd__clkbuf_4 _15200_ (.A(_07468_),
    .X(_07814_));
 sky130_fd_sc_hd__nor2_1 _15201_ (.A(_07814_),
    .B(_07685_),
    .Y(_07815_));
 sky130_fd_sc_hd__and2_1 _15202_ (.A(_07455_),
    .B(_07641_),
    .X(_07816_));
 sky130_fd_sc_hd__clkbuf_4 _15203_ (.A(_07816_),
    .X(_07817_));
 sky130_fd_sc_hd__nand2_1 _15204_ (.A(_07453_),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .Y(_07818_));
 sky130_fd_sc_hd__and2_1 _15205_ (.A(_07101_),
    .B(_07220_),
    .X(_07819_));
 sky130_fd_sc_hd__a21o_1 _15206_ (.A1(_07689_),
    .A2(_07690_),
    .B1(_07819_),
    .X(_07820_));
 sky130_fd_sc_hd__or3_1 _15207_ (.A(_07217_),
    .B(_07221_),
    .C(_07687_),
    .X(_07821_));
 sky130_fd_sc_hd__inv_2 _15208_ (.A(_07694_),
    .Y(_07822_));
 sky130_fd_sc_hd__a31o_1 _15209_ (.A1(_04933_),
    .A2(_07820_),
    .A3(_07821_),
    .B1(_07822_),
    .X(_07823_));
 sky130_fd_sc_hd__a21o_2 _15210_ (.A1(_07818_),
    .A2(_07823_),
    .B1(_07519_),
    .X(_07824_));
 sky130_fd_sc_hd__or4_1 _15211_ (.A(_07470_),
    .B(_07471_),
    .C(_07817_),
    .D(_07824_),
    .X(_07825_));
 sky130_fd_sc_hd__buf_4 _15212_ (.A(_07470_),
    .X(_07826_));
 sky130_fd_sc_hd__clkbuf_4 _15213_ (.A(_07824_),
    .X(_07827_));
 sky130_fd_sc_hd__o22ai_1 _15214_ (.A1(_07826_),
    .A2(_07817_),
    .B1(_07827_),
    .B2(_07471_),
    .Y(_07828_));
 sky130_fd_sc_hd__nand2_1 _15215_ (.A(_07825_),
    .B(_07828_),
    .Y(_07829_));
 sky130_fd_sc_hd__xnor2_1 _15216_ (.A(_07815_),
    .B(_07829_),
    .Y(_07830_));
 sky130_fd_sc_hd__nor2_1 _15217_ (.A(_03795_),
    .B(\rbzero.wall_tracer.stepDistY[2] ),
    .Y(_07831_));
 sky130_fd_sc_hd__inv_2 _15218_ (.A(_07831_),
    .Y(_07832_));
 sky130_fd_sc_hd__and2_1 _15219_ (.A(_04937_),
    .B(\rbzero.wall_tracer.stepDistX[2] ),
    .X(_07833_));
 sky130_fd_sc_hd__a31oi_4 _15220_ (.A1(_04928_),
    .A2(_07832_),
    .A3(_07651_),
    .B1(_07833_),
    .Y(_07834_));
 sky130_fd_sc_hd__buf_4 _15221_ (.A(_07646_),
    .X(_07835_));
 sky130_fd_sc_hd__or4_1 _15222_ (.A(_07834_),
    .B(_07835_),
    .C(_07663_),
    .D(_07680_),
    .X(_07836_));
 sky130_fd_sc_hd__a31o_2 _15223_ (.A1(_04929_),
    .A2(_07832_),
    .A3(_07651_),
    .B1(_07833_),
    .X(_07837_));
 sky130_fd_sc_hd__a21o_4 _15224_ (.A1(\rbzero.debug_overlay.playerX[-9] ),
    .A2(_04937_),
    .B1(_07643_),
    .X(_07838_));
 sky130_fd_sc_hd__a2bb2o_1 _15225_ (.A1_N(_07663_),
    .A2_N(_07680_),
    .B1(_07837_),
    .B2(_07838_),
    .X(_07839_));
 sky130_fd_sc_hd__nor2_2 _15226_ (.A(_07686_),
    .B(_07695_),
    .Y(_07840_));
 sky130_fd_sc_hd__or2_1 _15227_ (.A(_04935_),
    .B(_07664_),
    .X(_07841_));
 sky130_fd_sc_hd__buf_2 _15228_ (.A(_07841_),
    .X(_07842_));
 sky130_fd_sc_hd__buf_4 _15229_ (.A(_07842_),
    .X(_07843_));
 sky130_fd_sc_hd__nor2_1 _15230_ (.A(_07840_),
    .B(_07843_),
    .Y(_07844_));
 sky130_fd_sc_hd__nand3_1 _15231_ (.A(_07836_),
    .B(_07839_),
    .C(_07844_),
    .Y(_07845_));
 sky130_fd_sc_hd__a21o_1 _15232_ (.A1(_07836_),
    .A2(_07839_),
    .B1(_07844_),
    .X(_07846_));
 sky130_fd_sc_hd__clkbuf_4 _15233_ (.A(_07664_),
    .X(_07847_));
 sky130_fd_sc_hd__nand2_1 _15234_ (.A(_07647_),
    .B(_07653_),
    .Y(_07848_));
 sky130_fd_sc_hd__o31ai_1 _15235_ (.A1(_07663_),
    .A2(_07847_),
    .A3(_07654_),
    .B1(_07848_),
    .Y(_07849_));
 sky130_fd_sc_hd__nand3_1 _15236_ (.A(_07845_),
    .B(_07846_),
    .C(_07849_),
    .Y(_07850_));
 sky130_fd_sc_hd__a21o_1 _15237_ (.A1(_07845_),
    .A2(_07846_),
    .B1(_07849_),
    .X(_07851_));
 sky130_fd_sc_hd__nand3_1 _15238_ (.A(_07830_),
    .B(_07850_),
    .C(_07851_),
    .Y(_07852_));
 sky130_fd_sc_hd__a21o_1 _15239_ (.A1(_07850_),
    .A2(_07851_),
    .B1(_07830_),
    .X(_07853_));
 sky130_fd_sc_hd__nor2_1 _15240_ (.A(_07666_),
    .B(_07682_),
    .Y(_07854_));
 sky130_fd_sc_hd__a21o_1 _15241_ (.A1(_07683_),
    .A2(_07714_),
    .B1(_07854_),
    .X(_07855_));
 sky130_fd_sc_hd__nand3_1 _15242_ (.A(_07852_),
    .B(_07853_),
    .C(_07855_),
    .Y(_07856_));
 sky130_fd_sc_hd__a21o_1 _15243_ (.A1(_07852_),
    .A2(_07853_),
    .B1(_07855_),
    .X(_07857_));
 sky130_fd_sc_hd__clkbuf_4 _15244_ (.A(_07751_),
    .X(_07858_));
 sky130_fd_sc_hd__o31ai_2 _15245_ (.A1(_07469_),
    .A2(_07858_),
    .A3(_07750_),
    .B1(_07749_),
    .Y(_07859_));
 sky130_fd_sc_hd__inv_2 _15246_ (.A(_07713_),
    .Y(_07860_));
 sky130_fd_sc_hd__o21ba_1 _15247_ (.A1(_07700_),
    .A2(_07860_),
    .B1_N(_07699_),
    .X(_07861_));
 sky130_fd_sc_hd__nor2_1 _15248_ (.A(_07400_),
    .B(_07712_),
    .Y(_07862_));
 sky130_fd_sc_hd__o22a_1 _15249_ (.A1(_07379_),
    .A2(_07712_),
    .B1(_07736_),
    .B2(_07400_),
    .X(_07863_));
 sky130_fd_sc_hd__a21o_1 _15250_ (.A1(_07748_),
    .A2(_07862_),
    .B1(_07863_),
    .X(_07864_));
 sky130_fd_sc_hd__or2_1 _15251_ (.A(_07742_),
    .B(_07751_),
    .X(_07865_));
 sky130_fd_sc_hd__xor2_1 _15252_ (.A(_07864_),
    .B(_07865_),
    .X(_07866_));
 sky130_fd_sc_hd__xnor2_1 _15253_ (.A(_07861_),
    .B(_07866_),
    .Y(_07867_));
 sky130_fd_sc_hd__xor2_1 _15254_ (.A(_07859_),
    .B(_07867_),
    .X(_07868_));
 sky130_fd_sc_hd__nand3_1 _15255_ (.A(_07856_),
    .B(_07857_),
    .C(_07868_),
    .Y(_07869_));
 sky130_fd_sc_hd__a21o_1 _15256_ (.A1(_07856_),
    .A2(_07857_),
    .B1(_07868_),
    .X(_07870_));
 sky130_fd_sc_hd__nor2_1 _15257_ (.A(_07715_),
    .B(_07740_),
    .Y(_07871_));
 sky130_fd_sc_hd__a21o_1 _15258_ (.A1(_07741_),
    .A2(_07755_),
    .B1(_07871_),
    .X(_07872_));
 sky130_fd_sc_hd__nand3_1 _15259_ (.A(_07869_),
    .B(_07870_),
    .C(_07872_),
    .Y(_07873_));
 sky130_fd_sc_hd__a21o_1 _15260_ (.A1(_07869_),
    .A2(_07870_),
    .B1(_07872_),
    .X(_07874_));
 sky130_fd_sc_hd__a21o_1 _15261_ (.A1(_07798_),
    .A2(_07808_),
    .B1(_07807_),
    .X(_07875_));
 sky130_fd_sc_hd__nand2_1 _15262_ (.A(_07747_),
    .B(_07753_),
    .Y(_07876_));
 sky130_fd_sc_hd__or2b_1 _15263_ (.A(_07746_),
    .B_N(_07754_),
    .X(_07877_));
 sky130_fd_sc_hd__clkbuf_4 _15264_ (.A(_07792_),
    .X(_07878_));
 sky130_fd_sc_hd__and2_1 _15265_ (.A(_07571_),
    .B(_07572_),
    .X(_07879_));
 sky130_fd_sc_hd__clkbuf_4 _15266_ (.A(_07879_),
    .X(_07880_));
 sky130_fd_sc_hd__or4_1 _15267_ (.A(_07485_),
    .B(_07591_),
    .C(_07790_),
    .D(_07880_),
    .X(_07881_));
 sky130_fd_sc_hd__nand2_2 _15268_ (.A(_07571_),
    .B(_07572_),
    .Y(_07882_));
 sky130_fd_sc_hd__a22o_1 _15269_ (.A1(_07554_),
    .A2(_07793_),
    .B1(_07520_),
    .B2(_07882_),
    .X(_07883_));
 sky130_fd_sc_hd__nand2_1 _15270_ (.A(_07881_),
    .B(_07883_),
    .Y(_07884_));
 sky130_fd_sc_hd__or3_1 _15271_ (.A(_07878_),
    .B(_07598_),
    .C(_07884_),
    .X(_07885_));
 sky130_fd_sc_hd__clkbuf_4 _15272_ (.A(_07598_),
    .X(_07886_));
 sky130_fd_sc_hd__o21ai_1 _15273_ (.A1(_07878_),
    .A2(_07886_),
    .B1(_07884_),
    .Y(_07887_));
 sky130_fd_sc_hd__and2_1 _15274_ (.A(_07885_),
    .B(_07887_),
    .X(_07888_));
 sky130_fd_sc_hd__or4_1 _15275_ (.A(_07355_),
    .B(_07387_),
    .C(_07552_),
    .D(_07550_),
    .X(_07889_));
 sky130_fd_sc_hd__buf_2 _15276_ (.A(_07552_),
    .X(_07890_));
 sky130_fd_sc_hd__o22ai_1 _15277_ (.A1(_07469_),
    .A2(_07890_),
    .B1(_07800_),
    .B2(_07388_),
    .Y(_07891_));
 sky130_fd_sc_hd__nand2_1 _15278_ (.A(_07889_),
    .B(_07891_),
    .Y(_07892_));
 sky130_fd_sc_hd__or2_1 _15279_ (.A(_07424_),
    .B(_07567_),
    .X(_07893_));
 sky130_fd_sc_hd__xnor2_1 _15280_ (.A(_07892_),
    .B(_07893_),
    .Y(_07894_));
 sky130_fd_sc_hd__o31a_1 _15281_ (.A1(_07485_),
    .A2(_07805_),
    .A3(_07802_),
    .B1(_07799_),
    .X(_07895_));
 sky130_fd_sc_hd__nor2_1 _15282_ (.A(_07894_),
    .B(_07895_),
    .Y(_07896_));
 sky130_fd_sc_hd__nand2_1 _15283_ (.A(_07894_),
    .B(_07895_),
    .Y(_07897_));
 sky130_fd_sc_hd__and2b_1 _15284_ (.A_N(_07896_),
    .B(_07897_),
    .X(_07898_));
 sky130_fd_sc_hd__xnor2_1 _15285_ (.A(_07888_),
    .B(_07898_),
    .Y(_07899_));
 sky130_fd_sc_hd__a21o_1 _15286_ (.A1(_07876_),
    .A2(_07877_),
    .B1(_07899_),
    .X(_07900_));
 sky130_fd_sc_hd__nand3_1 _15287_ (.A(_07876_),
    .B(_07877_),
    .C(_07899_),
    .Y(_07901_));
 sky130_fd_sc_hd__nand2_1 _15288_ (.A(_07900_),
    .B(_07901_),
    .Y(_07902_));
 sky130_fd_sc_hd__xnor2_1 _15289_ (.A(_07875_),
    .B(_07902_),
    .Y(_07903_));
 sky130_fd_sc_hd__nand3_1 _15290_ (.A(_07873_),
    .B(_07874_),
    .C(_07903_),
    .Y(_07904_));
 sky130_fd_sc_hd__a21o_1 _15291_ (.A1(_07873_),
    .A2(_07874_),
    .B1(_07903_),
    .X(_07905_));
 sky130_fd_sc_hd__o211ai_1 _15292_ (.A1(_07782_),
    .A2(_07813_),
    .B1(_07904_),
    .C1(_07905_),
    .Y(_07906_));
 sky130_fd_sc_hd__a211o_1 _15293_ (.A1(_07904_),
    .A2(_07905_),
    .B1(_07782_),
    .C1(_07813_),
    .X(_07907_));
 sky130_fd_sc_hd__or2b_1 _15294_ (.A(_07810_),
    .B_N(_07787_),
    .X(_07908_));
 sky130_fd_sc_hd__or2b_1 _15295_ (.A(_07811_),
    .B_N(_07784_),
    .X(_07909_));
 sky130_fd_sc_hd__or4b_1 _15296_ (.A(_07517_),
    .B(_07529_),
    .C(_07620_),
    .D_N(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_07910_));
 sky130_fd_sc_hd__inv_2 _15297_ (.A(_07910_),
    .Y(_07911_));
 sky130_fd_sc_hd__o22a_1 _15298_ (.A1(_07616_),
    .A2(_07617_),
    .B1(_07621_),
    .B2(_07788_),
    .X(_07912_));
 sky130_fd_sc_hd__nor2_1 _15299_ (.A(_07911_),
    .B(_07912_),
    .Y(_07913_));
 sky130_fd_sc_hd__nand2_4 _15300_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_03795_),
    .Y(_07914_));
 sky130_fd_sc_hd__or2_1 _15301_ (.A(_04937_),
    .B(_07914_),
    .X(_07915_));
 sky130_fd_sc_hd__buf_2 _15302_ (.A(_07915_),
    .X(_07916_));
 sky130_fd_sc_hd__nor2_1 _15303_ (.A(_07602_),
    .B(_07916_),
    .Y(_07917_));
 sky130_fd_sc_hd__xnor2_1 _15304_ (.A(_07913_),
    .B(_07917_),
    .Y(_07918_));
 sky130_fd_sc_hd__and3_1 _15305_ (.A(_07791_),
    .B(_07796_),
    .C(_07918_),
    .X(_07919_));
 sky130_fd_sc_hd__a21oi_1 _15306_ (.A1(_07791_),
    .A2(_07796_),
    .B1(_07918_),
    .Y(_07920_));
 sky130_fd_sc_hd__or2_1 _15307_ (.A(_07919_),
    .B(_07920_),
    .X(_07921_));
 sky130_fd_sc_hd__and2b_1 _15308_ (.A_N(_07623_),
    .B(_07628_),
    .X(_07922_));
 sky130_fd_sc_hd__xnor2_1 _15309_ (.A(_07921_),
    .B(_07922_),
    .Y(_07923_));
 sky130_fd_sc_hd__a21oi_1 _15310_ (.A1(_07908_),
    .A2(_07909_),
    .B1(_07923_),
    .Y(_07924_));
 sky130_fd_sc_hd__and3_1 _15311_ (.A(_07908_),
    .B(_07909_),
    .C(_07923_),
    .X(_07925_));
 sky130_fd_sc_hd__nor2_1 _15312_ (.A(_07924_),
    .B(_07925_),
    .Y(_07926_));
 sky130_fd_sc_hd__xnor2_1 _15313_ (.A(_07637_),
    .B(_07926_),
    .Y(_07927_));
 sky130_fd_sc_hd__nand3_1 _15314_ (.A(_07906_),
    .B(_07907_),
    .C(_07927_),
    .Y(_07928_));
 sky130_fd_sc_hd__a21o_1 _15315_ (.A1(_07906_),
    .A2(_07907_),
    .B1(_07927_),
    .X(_07929_));
 sky130_fd_sc_hd__nand2_1 _15316_ (.A(_07928_),
    .B(_07929_),
    .Y(_07930_));
 sky130_fd_sc_hd__xnor2_1 _15317_ (.A(_07783_),
    .B(_07812_),
    .Y(_07931_));
 sky130_fd_sc_hd__xnor2_1 _15318_ (.A(_07773_),
    .B(_07779_),
    .Y(_07932_));
 sky130_fd_sc_hd__xnor2_1 _15319_ (.A(_07764_),
    .B(_07770_),
    .Y(_07933_));
 sky130_fd_sc_hd__a2bb2o_1 _15320_ (.A1_N(_07760_),
    .A2_N(_07664_),
    .B1(_07759_),
    .B2(_07761_),
    .X(_07934_));
 sky130_fd_sc_hd__a211o_1 _15321_ (.A1(_07439_),
    .A2(_07440_),
    .B1(_07441_),
    .C1(_07645_),
    .X(_07935_));
 sky130_fd_sc_hd__nand2_2 _15322_ (.A(_07730_),
    .B(_07732_),
    .Y(_07936_));
 sky130_fd_sc_hd__nor2_1 _15323_ (.A(_07936_),
    .B(_07718_),
    .Y(_07937_));
 sky130_fd_sc_hd__xnor2_1 _15324_ (.A(_07935_),
    .B(_07937_),
    .Y(_07938_));
 sky130_fd_sc_hd__nor2_1 _15325_ (.A(_07664_),
    .B(_07709_),
    .Y(_07939_));
 sky130_fd_sc_hd__or3_1 _15326_ (.A(_07936_),
    .B(_07718_),
    .C(_07935_),
    .X(_07940_));
 sky130_fd_sc_hd__a21bo_1 _15327_ (.A1(_07938_),
    .A2(_07939_),
    .B1_N(_07940_),
    .X(_07941_));
 sky130_fd_sc_hd__nand3_1 _15328_ (.A(_07762_),
    .B(_07934_),
    .C(_07941_),
    .Y(_07942_));
 sky130_fd_sc_hd__a21o_1 _15329_ (.A1(_07762_),
    .A2(_07934_),
    .B1(_07941_),
    .X(_07943_));
 sky130_fd_sc_hd__a2bb2o_1 _15330_ (.A1_N(_07468_),
    .A2_N(_07469_),
    .B1(_07456_),
    .B2(_07473_),
    .X(_07944_));
 sky130_fd_sc_hd__nand4_1 _15331_ (.A(_07474_),
    .B(_07942_),
    .C(_07943_),
    .D(_07944_),
    .Y(_07945_));
 sky130_fd_sc_hd__and2_1 _15332_ (.A(_07942_),
    .B(_07945_),
    .X(_07946_));
 sky130_fd_sc_hd__xor2_1 _15333_ (.A(_07933_),
    .B(_07946_),
    .X(_07947_));
 sky130_fd_sc_hd__xor2_1 _15334_ (.A(_07488_),
    .B(_07489_),
    .X(_07948_));
 sky130_fd_sc_hd__nor2_1 _15335_ (.A(_07933_),
    .B(_07946_),
    .Y(_07949_));
 sky130_fd_sc_hd__a21oi_1 _15336_ (.A1(_07947_),
    .A2(_07948_),
    .B1(_07949_),
    .Y(_07950_));
 sky130_fd_sc_hd__xor2_1 _15337_ (.A(_07932_),
    .B(_07950_),
    .X(_07951_));
 sky130_fd_sc_hd__xnor2_1 _15338_ (.A(_07614_),
    .B(_07590_),
    .Y(_07952_));
 sky130_fd_sc_hd__nor2_1 _15339_ (.A(_07932_),
    .B(_07950_),
    .Y(_07953_));
 sky130_fd_sc_hd__a21oi_1 _15340_ (.A1(_07951_),
    .A2(_07952_),
    .B1(_07953_),
    .Y(_07954_));
 sky130_fd_sc_hd__xor2_1 _15341_ (.A(_07931_),
    .B(_07954_),
    .X(_07955_));
 sky130_fd_sc_hd__and3_1 _15342_ (.A(_07588_),
    .B(_07615_),
    .C(_07639_),
    .X(_07956_));
 sky130_fd_sc_hd__nor2_1 _15343_ (.A(_07640_),
    .B(_07956_),
    .Y(_07957_));
 sky130_fd_sc_hd__nor2_1 _15344_ (.A(_07931_),
    .B(_07954_),
    .Y(_07958_));
 sky130_fd_sc_hd__a21o_1 _15345_ (.A1(_07955_),
    .A2(_07957_),
    .B1(_07958_),
    .X(_07959_));
 sky130_fd_sc_hd__xnor2_1 _15346_ (.A(_07930_),
    .B(_07959_),
    .Y(_07960_));
 sky130_fd_sc_hd__xnor2_2 _15347_ (.A(_07640_),
    .B(_07960_),
    .Y(_07961_));
 sky130_fd_sc_hd__and2b_1 _15348_ (.A_N(_07613_),
    .B(_07612_),
    .X(_07962_));
 sky130_fd_sc_hd__xnor2_1 _15349_ (.A(_07604_),
    .B(_07962_),
    .Y(_07963_));
 sky130_fd_sc_hd__o31a_2 _15350_ (.A1(_04936_),
    .A2(_07392_),
    .A3(_07393_),
    .B1(_07397_),
    .X(_07964_));
 sky130_fd_sc_hd__a2bb2o_1 _15351_ (.A1_N(_07378_),
    .A2_N(_07423_),
    .B1(_07554_),
    .B2(_07964_),
    .X(_07965_));
 sky130_fd_sc_hd__nor2_1 _15352_ (.A(_07416_),
    .B(_07575_),
    .Y(_07966_));
 sky130_fd_sc_hd__nor4_1 _15353_ (.A(_07378_),
    .B(_07399_),
    .C(_07423_),
    .D(_07485_),
    .Y(_07967_));
 sky130_fd_sc_hd__a21o_1 _15354_ (.A1(_07965_),
    .A2(_07966_),
    .B1(_07967_),
    .X(_07968_));
 sky130_fd_sc_hd__or2_1 _15355_ (.A(_07435_),
    .B(_07355_),
    .X(_07969_));
 sky130_fd_sc_hd__nand2_2 _15356_ (.A(_04928_),
    .B(_07698_),
    .Y(_07970_));
 sky130_fd_sc_hd__clkbuf_4 _15357_ (.A(_07970_),
    .X(_07971_));
 sky130_fd_sc_hd__or2_1 _15358_ (.A(_07670_),
    .B(_07971_),
    .X(_07972_));
 sky130_fd_sc_hd__xnor2_2 _15359_ (.A(_07969_),
    .B(_07972_),
    .Y(_07973_));
 sky130_fd_sc_hd__or2_1 _15360_ (.A(_07969_),
    .B(_07972_),
    .X(_07974_));
 sky130_fd_sc_hd__o31a_1 _15361_ (.A1(_07468_),
    .A2(_07388_),
    .A3(_07973_),
    .B1(_07974_),
    .X(_07975_));
 sky130_fd_sc_hd__nand2_1 _15362_ (.A(_07487_),
    .B(_07477_),
    .Y(_07976_));
 sky130_fd_sc_hd__xnor2_1 _15363_ (.A(_07976_),
    .B(_07486_),
    .Y(_07977_));
 sky130_fd_sc_hd__xnor2_1 _15364_ (.A(_07975_),
    .B(_07977_),
    .Y(_07978_));
 sky130_fd_sc_hd__or2b_1 _15365_ (.A(_07975_),
    .B_N(_07977_),
    .X(_07979_));
 sky130_fd_sc_hd__a21bo_1 _15366_ (.A1(_07968_),
    .A2(_07978_),
    .B1_N(_07979_),
    .X(_07980_));
 sky130_fd_sc_hd__or2b_1 _15367_ (.A(_07963_),
    .B_N(_07980_),
    .X(_07981_));
 sky130_fd_sc_hd__xor2_1 _15368_ (.A(_07980_),
    .B(_07963_),
    .X(_07982_));
 sky130_fd_sc_hd__a21oi_1 _15369_ (.A1(_07606_),
    .A2(_07608_),
    .B1(_07609_),
    .Y(_07983_));
 sky130_fd_sc_hd__nand2_1 _15370_ (.A(_04935_),
    .B(\rbzero.wall_tracer.stepDistX[-11] ),
    .Y(_07984_));
 sky130_fd_sc_hd__and2_1 _15371_ (.A(_07529_),
    .B(_07984_),
    .X(_07985_));
 sky130_fd_sc_hd__buf_2 _15372_ (.A(_07985_),
    .X(_07986_));
 sky130_fd_sc_hd__or4_1 _15373_ (.A(_07508_),
    .B(_07542_),
    .C(_07549_),
    .D(_07593_),
    .X(_07987_));
 sky130_fd_sc_hd__o22ai_1 _15374_ (.A1(_07508_),
    .A2(_07542_),
    .B1(_07550_),
    .B2(_07593_),
    .Y(_07988_));
 sky130_fd_sc_hd__nand2_1 _15375_ (.A(_07987_),
    .B(_07988_),
    .Y(_07989_));
 sky130_fd_sc_hd__o31a_1 _15376_ (.A1(_07567_),
    .A2(_07986_),
    .A3(_07989_),
    .B1(_07987_),
    .X(_07990_));
 sky130_fd_sc_hd__or2_1 _15377_ (.A(_07501_),
    .B(_07986_),
    .X(_07991_));
 sky130_fd_sc_hd__or3_1 _15378_ (.A(_07509_),
    .B(_07633_),
    .C(_07991_),
    .X(_07992_));
 sky130_fd_sc_hd__o21ai_1 _15379_ (.A1(_07509_),
    .A2(_07633_),
    .B1(_07991_),
    .Y(_07993_));
 sky130_fd_sc_hd__and2_1 _15380_ (.A(_07992_),
    .B(_07993_),
    .X(_07994_));
 sky130_fd_sc_hd__nor2_1 _15381_ (.A(_07610_),
    .B(_07983_),
    .Y(_07995_));
 sky130_fd_sc_hd__xnor2_1 _15382_ (.A(_07995_),
    .B(_07990_),
    .Y(_07996_));
 sky130_fd_sc_hd__nand2_1 _15383_ (.A(_07994_),
    .B(_07996_),
    .Y(_07997_));
 sky130_fd_sc_hd__o31ai_1 _15384_ (.A1(_07610_),
    .A2(_07983_),
    .A3(_07990_),
    .B1(_07997_),
    .Y(_07998_));
 sky130_fd_sc_hd__or2b_1 _15385_ (.A(_07982_),
    .B_N(_07998_),
    .X(_07999_));
 sky130_fd_sc_hd__and2_1 _15386_ (.A(_07622_),
    .B(_07635_),
    .X(_08000_));
 sky130_fd_sc_hd__or2_1 _15387_ (.A(_07636_),
    .B(_08000_),
    .X(_08001_));
 sky130_fd_sc_hd__a21oi_2 _15388_ (.A1(_07981_),
    .A2(_07999_),
    .B1(_08001_),
    .Y(_08002_));
 sky130_fd_sc_hd__xnor2_1 _15389_ (.A(_07955_),
    .B(_07957_),
    .Y(_08003_));
 sky130_fd_sc_hd__xnor2_1 _15390_ (.A(_07951_),
    .B(_07952_),
    .Y(_08004_));
 sky130_fd_sc_hd__xnor2_1 _15391_ (.A(_07947_),
    .B(_07948_),
    .Y(_08005_));
 sky130_fd_sc_hd__a22o_1 _15392_ (.A1(_07942_),
    .A2(_07943_),
    .B1(_07944_),
    .B2(_07474_),
    .X(_08006_));
 sky130_fd_sc_hd__xnor2_2 _15393_ (.A(_07938_),
    .B(_07939_),
    .Y(_08007_));
 sky130_fd_sc_hd__a211o_1 _15394_ (.A1(_07350_),
    .A2(_07353_),
    .B1(_07354_),
    .C1(_07644_),
    .X(_08008_));
 sky130_fd_sc_hd__a21oi_1 _15395_ (.A1(_07439_),
    .A2(_07440_),
    .B1(_07718_),
    .Y(_08009_));
 sky130_fd_sc_hd__xnor2_1 _15396_ (.A(_08008_),
    .B(_08009_),
    .Y(_08010_));
 sky130_fd_sc_hd__nor2_1 _15397_ (.A(_07842_),
    .B(_07936_),
    .Y(_08011_));
 sky130_fd_sc_hd__and2b_1 _15398_ (.A_N(_08008_),
    .B(_08009_),
    .X(_08012_));
 sky130_fd_sc_hd__a21oi_2 _15399_ (.A1(_08010_),
    .A2(_08011_),
    .B1(_08012_),
    .Y(_08013_));
 sky130_fd_sc_hd__xor2_2 _15400_ (.A(_08007_),
    .B(_08013_),
    .X(_08014_));
 sky130_fd_sc_hd__nor2_1 _15401_ (.A(_07468_),
    .B(_07388_),
    .Y(_08015_));
 sky130_fd_sc_hd__xnor2_2 _15402_ (.A(_07973_),
    .B(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__nor2_1 _15403_ (.A(_08007_),
    .B(_08013_),
    .Y(_08017_));
 sky130_fd_sc_hd__a21o_1 _15404_ (.A1(_08014_),
    .A2(_08016_),
    .B1(_08017_),
    .X(_08018_));
 sky130_fd_sc_hd__a21o_1 _15405_ (.A1(_07945_),
    .A2(_08006_),
    .B1(_08018_),
    .X(_08019_));
 sky130_fd_sc_hd__xor2_1 _15406_ (.A(_07968_),
    .B(_07978_),
    .X(_08020_));
 sky130_fd_sc_hd__nand3_1 _15407_ (.A(_07945_),
    .B(_08006_),
    .C(_08018_),
    .Y(_08021_));
 sky130_fd_sc_hd__a21boi_1 _15408_ (.A1(_08019_),
    .A2(_08020_),
    .B1_N(_08021_),
    .Y(_08022_));
 sky130_fd_sc_hd__xor2_1 _15409_ (.A(_08005_),
    .B(_08022_),
    .X(_08023_));
 sky130_fd_sc_hd__xnor2_1 _15410_ (.A(_07998_),
    .B(_07982_),
    .Y(_08024_));
 sky130_fd_sc_hd__nor2_1 _15411_ (.A(_08005_),
    .B(_08022_),
    .Y(_08025_));
 sky130_fd_sc_hd__a21oi_1 _15412_ (.A1(_08023_),
    .A2(_08024_),
    .B1(_08025_),
    .Y(_08026_));
 sky130_fd_sc_hd__xor2_1 _15413_ (.A(_08004_),
    .B(_08026_),
    .X(_08027_));
 sky130_fd_sc_hd__and3_1 _15414_ (.A(_07981_),
    .B(_07999_),
    .C(_08001_),
    .X(_08028_));
 sky130_fd_sc_hd__nor2_1 _15415_ (.A(_08002_),
    .B(_08028_),
    .Y(_08029_));
 sky130_fd_sc_hd__nor2_1 _15416_ (.A(_08004_),
    .B(_08026_),
    .Y(_08030_));
 sky130_fd_sc_hd__a21oi_1 _15417_ (.A1(_08027_),
    .A2(_08029_),
    .B1(_08030_),
    .Y(_08031_));
 sky130_fd_sc_hd__xor2_1 _15418_ (.A(_08003_),
    .B(_08031_),
    .X(_08032_));
 sky130_fd_sc_hd__nor2_1 _15419_ (.A(_08003_),
    .B(_08031_),
    .Y(_08033_));
 sky130_fd_sc_hd__a21oi_2 _15420_ (.A1(_08002_),
    .A2(_08032_),
    .B1(_08033_),
    .Y(_08034_));
 sky130_fd_sc_hd__xnor2_2 _15421_ (.A(_07961_),
    .B(_08034_),
    .Y(_08035_));
 sky130_fd_sc_hd__xnor2_1 _15422_ (.A(_08002_),
    .B(_08032_),
    .Y(_08036_));
 sky130_fd_sc_hd__nor2_1 _15423_ (.A(_07467_),
    .B(_07423_),
    .Y(_08037_));
 sky130_fd_sc_hd__or2_1 _15424_ (.A(_07435_),
    .B(_07387_),
    .X(_08038_));
 sky130_fd_sc_hd__nor2_1 _15425_ (.A(_07443_),
    .B(_07708_),
    .Y(_08039_));
 sky130_fd_sc_hd__xnor2_1 _15426_ (.A(_08038_),
    .B(_08039_),
    .Y(_08040_));
 sky130_fd_sc_hd__or3_1 _15427_ (.A(_07443_),
    .B(_07709_),
    .C(_08038_),
    .X(_08041_));
 sky130_fd_sc_hd__a21boi_1 _15428_ (.A1(_08037_),
    .A2(_08040_),
    .B1_N(_08041_),
    .Y(_08042_));
 sky130_fd_sc_hd__and2b_1 _15429_ (.A_N(_07967_),
    .B(_07965_),
    .X(_08043_));
 sky130_fd_sc_hd__xnor2_1 _15430_ (.A(_08043_),
    .B(_07966_),
    .Y(_08044_));
 sky130_fd_sc_hd__nand2_1 _15431_ (.A(_07964_),
    .B(_07554_),
    .Y(_08045_));
 sky130_fd_sc_hd__o31a_4 _15432_ (.A1(_04936_),
    .A2(_07362_),
    .A3(_07363_),
    .B1(_07376_),
    .X(_08046_));
 sky130_fd_sc_hd__nand2_1 _15433_ (.A(_08046_),
    .B(_07579_),
    .Y(_08047_));
 sky130_fd_sc_hd__or2_1 _15434_ (.A(_07416_),
    .B(_07508_),
    .X(_08048_));
 sky130_fd_sc_hd__o22a_1 _15435_ (.A1(_07377_),
    .A2(_07485_),
    .B1(_07574_),
    .B2(_07398_),
    .X(_08049_));
 sky130_fd_sc_hd__o22a_1 _15436_ (.A1(_08045_),
    .A2(_08047_),
    .B1(_08048_),
    .B2(_08049_),
    .X(_08050_));
 sky130_fd_sc_hd__xor2_1 _15437_ (.A(_08042_),
    .B(_08044_),
    .X(_08051_));
 sky130_fd_sc_hd__or2b_1 _15438_ (.A(_08050_),
    .B_N(_08051_),
    .X(_08052_));
 sky130_fd_sc_hd__o21ai_1 _15439_ (.A1(_08042_),
    .A2(_08044_),
    .B1(_08052_),
    .Y(_08053_));
 sky130_fd_sc_hd__or2_1 _15440_ (.A(_07994_),
    .B(_07996_),
    .X(_08054_));
 sky130_fd_sc_hd__and2_1 _15441_ (.A(_07997_),
    .B(_08054_),
    .X(_08055_));
 sky130_fd_sc_hd__xnor2_1 _15442_ (.A(_08053_),
    .B(_08055_),
    .Y(_08056_));
 sky130_fd_sc_hd__nor2_1 _15443_ (.A(_07567_),
    .B(_07986_),
    .Y(_08057_));
 sky130_fd_sc_hd__xor2_1 _15444_ (.A(_08057_),
    .B(_07989_),
    .X(_08058_));
 sky130_fd_sc_hd__a21boi_4 _15445_ (.A1(_04936_),
    .A2(\rbzero.wall_tracer.stepDistX[-12] ),
    .B1_N(_07633_),
    .Y(_08059_));
 sky130_fd_sc_hd__buf_2 _15446_ (.A(_08059_),
    .X(_08060_));
 sky130_fd_sc_hd__or2_1 _15447_ (.A(_07542_),
    .B(_07592_),
    .X(_08061_));
 sky130_fd_sc_hd__or2_1 _15448_ (.A(_07549_),
    .B(_07986_),
    .X(_08062_));
 sky130_fd_sc_hd__or4_1 _15449_ (.A(_07542_),
    .B(_07549_),
    .C(_07592_),
    .D(_07985_),
    .X(_08063_));
 sky130_fd_sc_hd__a21bo_1 _15450_ (.A1(_08061_),
    .A2(_08062_),
    .B1_N(_08063_),
    .X(_08064_));
 sky130_fd_sc_hd__o31a_1 _15451_ (.A1(_07567_),
    .A2(_08060_),
    .A3(_08064_),
    .B1(_08063_),
    .X(_08065_));
 sky130_fd_sc_hd__xnor2_1 _15452_ (.A(_08058_),
    .B(_08065_),
    .Y(_08066_));
 sky130_fd_sc_hd__clkbuf_4 _15453_ (.A(_07591_),
    .X(_08067_));
 sky130_fd_sc_hd__or2_1 _15454_ (.A(_08067_),
    .B(_08060_),
    .X(_08068_));
 sky130_fd_sc_hd__or2_1 _15455_ (.A(_08058_),
    .B(_08065_),
    .X(_08069_));
 sky130_fd_sc_hd__o21ai_1 _15456_ (.A1(_08066_),
    .A2(_08068_),
    .B1(_08069_),
    .Y(_08070_));
 sky130_fd_sc_hd__and2b_1 _15457_ (.A_N(_08056_),
    .B(_08070_),
    .X(_08071_));
 sky130_fd_sc_hd__a21oi_1 _15458_ (.A1(_08053_),
    .A2(_08055_),
    .B1(_08071_),
    .Y(_08072_));
 sky130_fd_sc_hd__nor2_1 _15459_ (.A(_07992_),
    .B(_08072_),
    .Y(_08073_));
 sky130_fd_sc_hd__xnor2_1 _15460_ (.A(_08027_),
    .B(_08029_),
    .Y(_08074_));
 sky130_fd_sc_hd__xnor2_1 _15461_ (.A(_08023_),
    .B(_08024_),
    .Y(_08075_));
 sky130_fd_sc_hd__and3_1 _15462_ (.A(_08021_),
    .B(_08019_),
    .C(_08020_),
    .X(_08076_));
 sky130_fd_sc_hd__a21oi_1 _15463_ (.A1(_08021_),
    .A2(_08019_),
    .B1(_08020_),
    .Y(_08077_));
 sky130_fd_sc_hd__or2_1 _15464_ (.A(_08076_),
    .B(_08077_),
    .X(_08078_));
 sky130_fd_sc_hd__xnor2_2 _15465_ (.A(_08014_),
    .B(_08016_),
    .Y(_08079_));
 sky130_fd_sc_hd__xor2_1 _15466_ (.A(_08037_),
    .B(_08040_),
    .X(_08080_));
 sky130_fd_sc_hd__xnor2_1 _15467_ (.A(_08010_),
    .B(_08011_),
    .Y(_08081_));
 sky130_fd_sc_hd__a211o_1 _15468_ (.A1(_07384_),
    .A2(_07385_),
    .B1(_07386_),
    .C1(_07645_),
    .X(_08082_));
 sky130_fd_sc_hd__or4_1 _15469_ (.A(_07260_),
    .B(_07408_),
    .C(_04935_),
    .D(_07350_),
    .X(_08083_));
 sky130_fd_sc_hd__xor2_1 _15470_ (.A(_08082_),
    .B(_08083_),
    .X(_08084_));
 sky130_fd_sc_hd__and2_1 _15471_ (.A(_07439_),
    .B(_07440_),
    .X(_08085_));
 sky130_fd_sc_hd__clkbuf_4 _15472_ (.A(_08085_),
    .X(_08086_));
 sky130_fd_sc_hd__nor2_1 _15473_ (.A(_08086_),
    .B(_07842_),
    .Y(_08087_));
 sky130_fd_sc_hd__nor2_1 _15474_ (.A(_08082_),
    .B(_08083_),
    .Y(_08088_));
 sky130_fd_sc_hd__a21o_1 _15475_ (.A1(_08084_),
    .A2(_08087_),
    .B1(_08088_),
    .X(_08089_));
 sky130_fd_sc_hd__xnor2_1 _15476_ (.A(_08081_),
    .B(_08089_),
    .Y(_08090_));
 sky130_fd_sc_hd__and2b_1 _15477_ (.A_N(_08081_),
    .B(_08089_),
    .X(_08091_));
 sky130_fd_sc_hd__a21o_1 _15478_ (.A1(_08080_),
    .A2(_08090_),
    .B1(_08091_),
    .X(_08092_));
 sky130_fd_sc_hd__xnor2_2 _15479_ (.A(_08079_),
    .B(_08092_),
    .Y(_08093_));
 sky130_fd_sc_hd__xnor2_1 _15480_ (.A(_08050_),
    .B(_08051_),
    .Y(_08094_));
 sky130_fd_sc_hd__and2b_1 _15481_ (.A_N(_08079_),
    .B(_08092_),
    .X(_08095_));
 sky130_fd_sc_hd__a21oi_1 _15482_ (.A1(_08093_),
    .A2(_08094_),
    .B1(_08095_),
    .Y(_08096_));
 sky130_fd_sc_hd__xor2_1 _15483_ (.A(_08078_),
    .B(_08096_),
    .X(_08097_));
 sky130_fd_sc_hd__xnor2_1 _15484_ (.A(_08070_),
    .B(_08056_),
    .Y(_08098_));
 sky130_fd_sc_hd__nor2_1 _15485_ (.A(_08078_),
    .B(_08096_),
    .Y(_08099_));
 sky130_fd_sc_hd__a21oi_1 _15486_ (.A1(_08097_),
    .A2(_08098_),
    .B1(_08099_),
    .Y(_08100_));
 sky130_fd_sc_hd__nand2_1 _15487_ (.A(_08075_),
    .B(_08100_),
    .Y(_08101_));
 sky130_fd_sc_hd__and2_1 _15488_ (.A(_07992_),
    .B(_08072_),
    .X(_08102_));
 sky130_fd_sc_hd__nor2_1 _15489_ (.A(_08073_),
    .B(_08102_),
    .Y(_08103_));
 sky130_fd_sc_hd__nor2_1 _15490_ (.A(_08075_),
    .B(_08100_),
    .Y(_08104_));
 sky130_fd_sc_hd__a21o_1 _15491_ (.A1(_08101_),
    .A2(_08103_),
    .B1(_08104_),
    .X(_08105_));
 sky130_fd_sc_hd__xnor2_1 _15492_ (.A(_08074_),
    .B(_08105_),
    .Y(_08106_));
 sky130_fd_sc_hd__or2b_1 _15493_ (.A(_08074_),
    .B_N(_08105_),
    .X(_08107_));
 sky130_fd_sc_hd__a21boi_1 _15494_ (.A1(_08073_),
    .A2(_08106_),
    .B1_N(_08107_),
    .Y(_08108_));
 sky130_fd_sc_hd__or2_1 _15495_ (.A(_08036_),
    .B(_08108_),
    .X(_08109_));
 sky130_fd_sc_hd__nand2_1 _15496_ (.A(_08035_),
    .B(_08109_),
    .Y(_08110_));
 sky130_fd_sc_hd__xor2_1 _15497_ (.A(_08036_),
    .B(_08108_),
    .X(_08111_));
 sky130_fd_sc_hd__xor2_1 _15498_ (.A(_08073_),
    .B(_08106_),
    .X(_08112_));
 sky130_fd_sc_hd__and2b_1 _15499_ (.A_N(_08104_),
    .B(_08101_),
    .X(_08113_));
 sky130_fd_sc_hd__xnor2_1 _15500_ (.A(_08113_),
    .B(_08103_),
    .Y(_08114_));
 sky130_fd_sc_hd__xnor2_1 _15501_ (.A(_08097_),
    .B(_08098_),
    .Y(_08115_));
 sky130_fd_sc_hd__xnor2_2 _15502_ (.A(_08093_),
    .B(_08094_),
    .Y(_08116_));
 sky130_fd_sc_hd__nor2_1 _15503_ (.A(_07416_),
    .B(_07593_),
    .Y(_08117_));
 sky130_fd_sc_hd__nor4_1 _15504_ (.A(_07378_),
    .B(_07399_),
    .C(_07508_),
    .D(_07575_),
    .Y(_08118_));
 sky130_fd_sc_hd__o22a_1 _15505_ (.A1(_07399_),
    .A2(_07508_),
    .B1(_07575_),
    .B2(_07378_),
    .X(_08119_));
 sky130_fd_sc_hd__nor2_1 _15506_ (.A(_08118_),
    .B(_08119_),
    .Y(_08120_));
 sky130_fd_sc_hd__a21o_1 _15507_ (.A1(_08117_),
    .A2(_08120_),
    .B1(_08118_),
    .X(_08121_));
 sky130_fd_sc_hd__nor2_1 _15508_ (.A(_07467_),
    .B(_07485_),
    .Y(_08122_));
 sky130_fd_sc_hd__nor2_2 _15509_ (.A(_04936_),
    .B(_07733_),
    .Y(_08123_));
 sky130_fd_sc_hd__a2bb2o_1 _15510_ (.A1_N(_07435_),
    .A2_N(_07423_),
    .B1(_08123_),
    .B2(_07698_),
    .X(_08124_));
 sky130_fd_sc_hd__or4_1 _15511_ (.A(_07435_),
    .B(_07423_),
    .C(_07970_),
    .D(_07936_),
    .X(_08125_));
 sky130_fd_sc_hd__a21boi_1 _15512_ (.A1(_08122_),
    .A2(_08124_),
    .B1_N(_08125_),
    .Y(_08126_));
 sky130_fd_sc_hd__o21ba_1 _15513_ (.A1(_08045_),
    .A2(_08047_),
    .B1_N(_08049_),
    .X(_08127_));
 sky130_fd_sc_hd__xor2_1 _15514_ (.A(_08048_),
    .B(_08127_),
    .X(_08128_));
 sky130_fd_sc_hd__xor2_1 _15515_ (.A(_08126_),
    .B(_08128_),
    .X(_08129_));
 sky130_fd_sc_hd__xor2_1 _15516_ (.A(_08121_),
    .B(_08129_),
    .X(_08130_));
 sky130_fd_sc_hd__xnor2_1 _15517_ (.A(_08080_),
    .B(_08090_),
    .Y(_08131_));
 sky130_fd_sc_hd__and2_1 _15518_ (.A(_08125_),
    .B(_08124_),
    .X(_08132_));
 sky130_fd_sc_hd__xor2_1 _15519_ (.A(_08122_),
    .B(_08132_),
    .X(_08133_));
 sky130_fd_sc_hd__xnor2_1 _15520_ (.A(_08084_),
    .B(_08087_),
    .Y(_08134_));
 sky130_fd_sc_hd__nand2_4 _15521_ (.A(_07350_),
    .B(_07353_),
    .Y(_08135_));
 sky130_fd_sc_hd__nor2_2 _15522_ (.A(_07466_),
    .B(_07664_),
    .Y(_08136_));
 sky130_fd_sc_hd__a211o_1 _15523_ (.A1(_07420_),
    .A2(_07421_),
    .B1(_07422_),
    .C1(_07645_),
    .X(_08137_));
 sky130_fd_sc_hd__or4_2 _15524_ (.A(_07260_),
    .B(_07408_),
    .C(_04935_),
    .D(_07384_),
    .X(_08138_));
 sky130_fd_sc_hd__xor2_2 _15525_ (.A(_08137_),
    .B(_08138_),
    .X(_08139_));
 sky130_fd_sc_hd__nor2_1 _15526_ (.A(_08137_),
    .B(_08138_),
    .Y(_08140_));
 sky130_fd_sc_hd__a31oi_2 _15527_ (.A1(_08135_),
    .A2(_08136_),
    .A3(_08139_),
    .B1(_08140_),
    .Y(_08141_));
 sky130_fd_sc_hd__xor2_1 _15528_ (.A(_08134_),
    .B(_08141_),
    .X(_08142_));
 sky130_fd_sc_hd__nor2_1 _15529_ (.A(_08134_),
    .B(_08141_),
    .Y(_08143_));
 sky130_fd_sc_hd__a21o_1 _15530_ (.A1(_08133_),
    .A2(_08142_),
    .B1(_08143_),
    .X(_08144_));
 sky130_fd_sc_hd__xnor2_1 _15531_ (.A(_08131_),
    .B(_08144_),
    .Y(_08145_));
 sky130_fd_sc_hd__and2b_1 _15532_ (.A_N(_08131_),
    .B(_08144_),
    .X(_08146_));
 sky130_fd_sc_hd__a21oi_2 _15533_ (.A1(_08130_),
    .A2(_08145_),
    .B1(_08146_),
    .Y(_08147_));
 sky130_fd_sc_hd__xor2_2 _15534_ (.A(_08116_),
    .B(_08147_),
    .X(_08148_));
 sky130_fd_sc_hd__nor2_1 _15535_ (.A(_08126_),
    .B(_08128_),
    .Y(_08149_));
 sky130_fd_sc_hd__a21o_1 _15536_ (.A1(_08121_),
    .A2(_08129_),
    .B1(_08149_),
    .X(_08150_));
 sky130_fd_sc_hd__xnor2_1 _15537_ (.A(_08066_),
    .B(_08068_),
    .Y(_08151_));
 sky130_fd_sc_hd__xor2_1 _15538_ (.A(_08150_),
    .B(_08151_),
    .X(_08152_));
 sky130_fd_sc_hd__nor2_1 _15539_ (.A(_07566_),
    .B(_08060_),
    .Y(_08153_));
 sky130_fd_sc_hd__xnor2_1 _15540_ (.A(_08153_),
    .B(_08064_),
    .Y(_08154_));
 sky130_fd_sc_hd__nor2_1 _15541_ (.A(_07552_),
    .B(_08059_),
    .Y(_08155_));
 sky130_fd_sc_hd__and2b_1 _15542_ (.A_N(_08062_),
    .B(_08155_),
    .X(_08156_));
 sky130_fd_sc_hd__and2_1 _15543_ (.A(_08154_),
    .B(_08156_),
    .X(_08157_));
 sky130_fd_sc_hd__xnor2_2 _15544_ (.A(_08152_),
    .B(_08157_),
    .Y(_08158_));
 sky130_fd_sc_hd__nor2_1 _15545_ (.A(_08116_),
    .B(_08147_),
    .Y(_08159_));
 sky130_fd_sc_hd__a21oi_1 _15546_ (.A1(_08148_),
    .A2(_08158_),
    .B1(_08159_),
    .Y(_08160_));
 sky130_fd_sc_hd__xnor2_1 _15547_ (.A(_08115_),
    .B(_08160_),
    .Y(_08161_));
 sky130_fd_sc_hd__or2b_1 _15548_ (.A(_08150_),
    .B_N(_08151_),
    .X(_08162_));
 sky130_fd_sc_hd__and2b_1 _15549_ (.A_N(_08151_),
    .B(_08150_),
    .X(_08163_));
 sky130_fd_sc_hd__a21oi_1 _15550_ (.A1(_08162_),
    .A2(_08157_),
    .B1(_08163_),
    .Y(_08164_));
 sky130_fd_sc_hd__or2_1 _15551_ (.A(_08115_),
    .B(_08160_),
    .X(_08165_));
 sky130_fd_sc_hd__o21a_1 _15552_ (.A1(_08161_),
    .A2(_08164_),
    .B1(_08165_),
    .X(_08166_));
 sky130_fd_sc_hd__nor2_1 _15553_ (.A(_08114_),
    .B(_08166_),
    .Y(_08167_));
 sky130_fd_sc_hd__and2_1 _15554_ (.A(_08112_),
    .B(_08167_),
    .X(_08168_));
 sky130_fd_sc_hd__nand2_1 _15555_ (.A(_08111_),
    .B(_08168_),
    .Y(_08169_));
 sky130_fd_sc_hd__or2_1 _15556_ (.A(_08111_),
    .B(_08168_),
    .X(_08170_));
 sky130_fd_sc_hd__and2_2 _15557_ (.A(_08169_),
    .B(_08170_),
    .X(_08171_));
 sky130_fd_sc_hd__xnor2_1 _15558_ (.A(_08114_),
    .B(_08166_),
    .Y(_08172_));
 sky130_fd_sc_hd__xnor2_1 _15559_ (.A(_08161_),
    .B(_08164_),
    .Y(_08173_));
 sky130_fd_sc_hd__nor2_1 _15560_ (.A(_07467_),
    .B(_07575_),
    .Y(_08174_));
 sky130_fd_sc_hd__a2bb2o_1 _15561_ (.A1_N(_08086_),
    .A2_N(_07970_),
    .B1(_07554_),
    .B2(_07697_),
    .X(_08175_));
 sky130_fd_sc_hd__or4_1 _15562_ (.A(_07435_),
    .B(_08086_),
    .C(_07484_),
    .D(_07970_),
    .X(_08176_));
 sky130_fd_sc_hd__a21boi_1 _15563_ (.A1(_08174_),
    .A2(_08175_),
    .B1_N(_08176_),
    .Y(_08177_));
 sky130_fd_sc_hd__xnor2_1 _15564_ (.A(_08117_),
    .B(_08120_),
    .Y(_08178_));
 sky130_fd_sc_hd__or2_1 _15565_ (.A(_08177_),
    .B(_08178_),
    .X(_08179_));
 sky130_fd_sc_hd__nor2_1 _15566_ (.A(_07416_),
    .B(_07986_),
    .Y(_08180_));
 sky130_fd_sc_hd__o22ai_1 _15567_ (.A1(_07378_),
    .A2(_07507_),
    .B1(_07592_),
    .B2(_07399_),
    .Y(_08181_));
 sky130_fd_sc_hd__or4_1 _15568_ (.A(_07377_),
    .B(_07398_),
    .C(_07507_),
    .D(_07592_),
    .X(_08182_));
 sky130_fd_sc_hd__a21bo_1 _15569_ (.A1(_08180_),
    .A2(_08181_),
    .B1_N(_08182_),
    .X(_08183_));
 sky130_fd_sc_hd__xor2_1 _15570_ (.A(_08177_),
    .B(_08178_),
    .X(_08184_));
 sky130_fd_sc_hd__nand2_1 _15571_ (.A(_08183_),
    .B(_08184_),
    .Y(_08185_));
 sky130_fd_sc_hd__nor2_1 _15572_ (.A(_08154_),
    .B(_08156_),
    .Y(_08186_));
 sky130_fd_sc_hd__or2_1 _15573_ (.A(_08157_),
    .B(_08186_),
    .X(_08187_));
 sky130_fd_sc_hd__a21oi_2 _15574_ (.A1(_08179_),
    .A2(_08185_),
    .B1(_08187_),
    .Y(_08188_));
 sky130_fd_sc_hd__xnor2_2 _15575_ (.A(_08148_),
    .B(_08158_),
    .Y(_08189_));
 sky130_fd_sc_hd__and3_1 _15576_ (.A(_08179_),
    .B(_08185_),
    .C(_08187_),
    .X(_08190_));
 sky130_fd_sc_hd__nor2_1 _15577_ (.A(_08188_),
    .B(_08190_),
    .Y(_08191_));
 sky130_fd_sc_hd__xnor2_1 _15578_ (.A(_08130_),
    .B(_08145_),
    .Y(_08192_));
 sky130_fd_sc_hd__xor2_1 _15579_ (.A(_08183_),
    .B(_08184_),
    .X(_08193_));
 sky130_fd_sc_hd__xnor2_1 _15580_ (.A(_08133_),
    .B(_08142_),
    .Y(_08194_));
 sky130_fd_sc_hd__and2_1 _15581_ (.A(_08176_),
    .B(_08175_),
    .X(_08195_));
 sky130_fd_sc_hd__xor2_2 _15582_ (.A(_08174_),
    .B(_08195_),
    .X(_08196_));
 sky130_fd_sc_hd__nand2_1 _15583_ (.A(_08135_),
    .B(_08136_),
    .Y(_08197_));
 sky130_fd_sc_hd__xor2_2 _15584_ (.A(_08139_),
    .B(_08197_),
    .X(_08198_));
 sky130_fd_sc_hd__a211o_1 _15585_ (.A1(_07481_),
    .A2(_07482_),
    .B1(_07483_),
    .C1(_07645_),
    .X(_08199_));
 sky130_fd_sc_hd__or4_2 _15586_ (.A(_07260_),
    .B(_07408_),
    .C(_07356_),
    .D(_07420_),
    .X(_08200_));
 sky130_fd_sc_hd__xor2_2 _15587_ (.A(_08199_),
    .B(_08200_),
    .X(_08201_));
 sky130_fd_sc_hd__and2_1 _15588_ (.A(_07384_),
    .B(_07385_),
    .X(_08202_));
 sky130_fd_sc_hd__nor2_1 _15589_ (.A(_08202_),
    .B(_07842_),
    .Y(_08203_));
 sky130_fd_sc_hd__nor2_1 _15590_ (.A(_08199_),
    .B(_08200_),
    .Y(_08204_));
 sky130_fd_sc_hd__a21oi_2 _15591_ (.A1(_08201_),
    .A2(_08203_),
    .B1(_08204_),
    .Y(_08205_));
 sky130_fd_sc_hd__xor2_2 _15592_ (.A(_08198_),
    .B(_08205_),
    .X(_08206_));
 sky130_fd_sc_hd__nor2_1 _15593_ (.A(_08198_),
    .B(_08205_),
    .Y(_08207_));
 sky130_fd_sc_hd__a21oi_1 _15594_ (.A1(_08196_),
    .A2(_08206_),
    .B1(_08207_),
    .Y(_08208_));
 sky130_fd_sc_hd__xor2_1 _15595_ (.A(_08194_),
    .B(_08208_),
    .X(_08209_));
 sky130_fd_sc_hd__nor2_1 _15596_ (.A(_08194_),
    .B(_08208_),
    .Y(_08210_));
 sky130_fd_sc_hd__a21o_1 _15597_ (.A1(_08193_),
    .A2(_08209_),
    .B1(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__xnor2_1 _15598_ (.A(_08192_),
    .B(_08211_),
    .Y(_08212_));
 sky130_fd_sc_hd__or2b_1 _15599_ (.A(_08192_),
    .B_N(_08211_),
    .X(_08213_));
 sky130_fd_sc_hd__a21boi_2 _15600_ (.A1(_08191_),
    .A2(_08212_),
    .B1_N(_08213_),
    .Y(_08214_));
 sky130_fd_sc_hd__xor2_2 _15601_ (.A(_08189_),
    .B(_08214_),
    .X(_08215_));
 sky130_fd_sc_hd__nor2_1 _15602_ (.A(_08189_),
    .B(_08214_),
    .Y(_08216_));
 sky130_fd_sc_hd__a21oi_1 _15603_ (.A1(_08188_),
    .A2(_08215_),
    .B1(_08216_),
    .Y(_08217_));
 sky130_fd_sc_hd__nor2_1 _15604_ (.A(_08173_),
    .B(_08217_),
    .Y(_08218_));
 sky130_fd_sc_hd__and2b_1 _15605_ (.A_N(_08172_),
    .B(_08218_),
    .X(_08219_));
 sky130_fd_sc_hd__and2_1 _15606_ (.A(_08173_),
    .B(_08217_),
    .X(_08220_));
 sky130_fd_sc_hd__nor2_2 _15607_ (.A(_08218_),
    .B(_08220_),
    .Y(_08221_));
 sky130_fd_sc_hd__and2_1 _15608_ (.A(_07350_),
    .B(_07353_),
    .X(_08222_));
 sky130_fd_sc_hd__clkbuf_4 _15609_ (.A(_08222_),
    .X(_08223_));
 sky130_fd_sc_hd__nor2_2 _15610_ (.A(_08223_),
    .B(_07971_),
    .Y(_08224_));
 sky130_fd_sc_hd__nand2_1 _15611_ (.A(_07697_),
    .B(_07579_),
    .Y(_08225_));
 sky130_fd_sc_hd__xnor2_2 _15612_ (.A(_08225_),
    .B(_08224_),
    .Y(_08226_));
 sky130_fd_sc_hd__nor2_1 _15613_ (.A(_07467_),
    .B(_07508_),
    .Y(_08227_));
 sky130_fd_sc_hd__a32oi_4 _15614_ (.A1(_07697_),
    .A2(_07579_),
    .A3(_08224_),
    .B1(_08226_),
    .B2(_08227_),
    .Y(_08228_));
 sky130_fd_sc_hd__and2_1 _15615_ (.A(_08182_),
    .B(_08181_),
    .X(_08229_));
 sky130_fd_sc_hd__xnor2_1 _15616_ (.A(_08180_),
    .B(_08229_),
    .Y(_08230_));
 sky130_fd_sc_hd__nor2_1 _15617_ (.A(_08228_),
    .B(_08230_),
    .Y(_08231_));
 sky130_fd_sc_hd__nor2_1 _15618_ (.A(_07416_),
    .B(_08059_),
    .Y(_08232_));
 sky130_fd_sc_hd__or2_1 _15619_ (.A(_07378_),
    .B(_07592_),
    .X(_08233_));
 sky130_fd_sc_hd__or2_1 _15620_ (.A(_07399_),
    .B(_07985_),
    .X(_08234_));
 sky130_fd_sc_hd__or4_1 _15621_ (.A(_07377_),
    .B(_07398_),
    .C(_07592_),
    .D(_07985_),
    .X(_08235_));
 sky130_fd_sc_hd__a21boi_1 _15622_ (.A1(_08233_),
    .A2(_08234_),
    .B1_N(_08235_),
    .Y(_08236_));
 sky130_fd_sc_hd__a21bo_1 _15623_ (.A1(_08232_),
    .A2(_08236_),
    .B1_N(_08235_),
    .X(_08237_));
 sky130_fd_sc_hd__xor2_1 _15624_ (.A(_08228_),
    .B(_08230_),
    .X(_08238_));
 sky130_fd_sc_hd__and2_1 _15625_ (.A(_08237_),
    .B(_08238_),
    .X(_08239_));
 sky130_fd_sc_hd__buf_4 _15626_ (.A(_07890_),
    .X(_08240_));
 sky130_fd_sc_hd__buf_4 _15627_ (.A(_07800_),
    .X(_08241_));
 sky130_fd_sc_hd__o22a_1 _15628_ (.A1(_08240_),
    .A2(_07986_),
    .B1(_08060_),
    .B2(_08241_),
    .X(_08242_));
 sky130_fd_sc_hd__nor2_1 _15629_ (.A(_08156_),
    .B(_08242_),
    .Y(_08243_));
 sky130_fd_sc_hd__o21a_1 _15630_ (.A1(_08231_),
    .A2(_08239_),
    .B1(_08243_),
    .X(_08244_));
 sky130_fd_sc_hd__xnor2_1 _15631_ (.A(_08191_),
    .B(_08212_),
    .Y(_08245_));
 sky130_fd_sc_hd__or3_1 _15632_ (.A(_08231_),
    .B(_08239_),
    .C(_08243_),
    .X(_08246_));
 sky130_fd_sc_hd__and2b_1 _15633_ (.A_N(_08244_),
    .B(_08246_),
    .X(_08247_));
 sky130_fd_sc_hd__xnor2_1 _15634_ (.A(_08193_),
    .B(_08209_),
    .Y(_08248_));
 sky130_fd_sc_hd__nand2_1 _15635_ (.A(_08196_),
    .B(_08206_),
    .Y(_08249_));
 sky130_fd_sc_hd__or2_1 _15636_ (.A(_08196_),
    .B(_08206_),
    .X(_08250_));
 sky130_fd_sc_hd__xor2_1 _15637_ (.A(_08227_),
    .B(_08226_),
    .X(_08251_));
 sky130_fd_sc_hd__xnor2_2 _15638_ (.A(_08201_),
    .B(_08203_),
    .Y(_08252_));
 sky130_fd_sc_hd__a211o_1 _15639_ (.A1(_07571_),
    .A2(_07572_),
    .B1(_07573_),
    .C1(_07645_),
    .X(_08253_));
 sky130_fd_sc_hd__or4_2 _15640_ (.A(_07260_),
    .B(_07453_),
    .C(_07356_),
    .D(_07481_),
    .X(_08254_));
 sky130_fd_sc_hd__xor2_1 _15641_ (.A(_08253_),
    .B(_08254_),
    .X(_08255_));
 sky130_fd_sc_hd__and2_2 _15642_ (.A(_07420_),
    .B(_07421_),
    .X(_08256_));
 sky130_fd_sc_hd__nor2_1 _15643_ (.A(_08256_),
    .B(_07842_),
    .Y(_08257_));
 sky130_fd_sc_hd__nor2_1 _15644_ (.A(_08253_),
    .B(_08254_),
    .Y(_08258_));
 sky130_fd_sc_hd__a21oi_1 _15645_ (.A1(_08255_),
    .A2(_08257_),
    .B1(_08258_),
    .Y(_08259_));
 sky130_fd_sc_hd__xor2_1 _15646_ (.A(_08252_),
    .B(_08259_),
    .X(_08260_));
 sky130_fd_sc_hd__nor2_1 _15647_ (.A(_08252_),
    .B(_08259_),
    .Y(_08261_));
 sky130_fd_sc_hd__a21o_1 _15648_ (.A1(_08251_),
    .A2(_08260_),
    .B1(_08261_),
    .X(_08262_));
 sky130_fd_sc_hd__xor2_1 _15649_ (.A(_08237_),
    .B(_08238_),
    .X(_08263_));
 sky130_fd_sc_hd__xnor2_1 _15650_ (.A(_08196_),
    .B(_08206_),
    .Y(_08264_));
 sky130_fd_sc_hd__xnor2_1 _15651_ (.A(_08264_),
    .B(_08262_),
    .Y(_08265_));
 sky130_fd_sc_hd__a32o_1 _15652_ (.A1(_08249_),
    .A2(_08250_),
    .A3(_08262_),
    .B1(_08263_),
    .B2(_08265_),
    .X(_08266_));
 sky130_fd_sc_hd__xnor2_1 _15653_ (.A(_08248_),
    .B(_08266_),
    .Y(_08267_));
 sky130_fd_sc_hd__or2b_1 _15654_ (.A(_08248_),
    .B_N(_08266_),
    .X(_08268_));
 sky130_fd_sc_hd__a21boi_1 _15655_ (.A1(_08247_),
    .A2(_08267_),
    .B1_N(_08268_),
    .Y(_08269_));
 sky130_fd_sc_hd__xor2_1 _15656_ (.A(_08245_),
    .B(_08269_),
    .X(_08270_));
 sky130_fd_sc_hd__xnor2_1 _15657_ (.A(_08244_),
    .B(_08270_),
    .Y(_08271_));
 sky130_fd_sc_hd__buf_4 _15658_ (.A(_07379_),
    .X(_08272_));
 sky130_fd_sc_hd__or2_1 _15659_ (.A(_07467_),
    .B(_07593_),
    .X(_08273_));
 sky130_fd_sc_hd__clkbuf_4 _15660_ (.A(_08202_),
    .X(_08274_));
 sky130_fd_sc_hd__or2_1 _15661_ (.A(_07435_),
    .B(_07507_),
    .X(_08275_));
 sky130_fd_sc_hd__o21a_1 _15662_ (.A1(_08274_),
    .A2(_07971_),
    .B1(_08275_),
    .X(_08276_));
 sky130_fd_sc_hd__or3_1 _15663_ (.A(_08274_),
    .B(_07971_),
    .C(_08275_),
    .X(_08277_));
 sky130_fd_sc_hd__o21a_1 _15664_ (.A1(_08273_),
    .A2(_08276_),
    .B1(_08277_),
    .X(_08278_));
 sky130_fd_sc_hd__xnor2_1 _15665_ (.A(_08232_),
    .B(_08236_),
    .Y(_08279_));
 sky130_fd_sc_hd__xnor2_1 _15666_ (.A(_08278_),
    .B(_08279_),
    .Y(_08280_));
 sky130_fd_sc_hd__or2_1 _15667_ (.A(_08278_),
    .B(_08279_),
    .X(_08281_));
 sky130_fd_sc_hd__o41a_1 _15668_ (.A1(_08272_),
    .A2(_08060_),
    .A3(_08234_),
    .A4(_08280_),
    .B1(_08281_),
    .X(_08282_));
 sky130_fd_sc_hd__and2b_1 _15669_ (.A_N(_08282_),
    .B(_08155_),
    .X(_08283_));
 sky130_fd_sc_hd__xnor2_1 _15670_ (.A(_08247_),
    .B(_08267_),
    .Y(_08284_));
 sky130_fd_sc_hd__and2b_1 _15671_ (.A_N(_08155_),
    .B(_08282_),
    .X(_08285_));
 sky130_fd_sc_hd__nor2_1 _15672_ (.A(_08283_),
    .B(_08285_),
    .Y(_08286_));
 sky130_fd_sc_hd__xnor2_1 _15673_ (.A(_08263_),
    .B(_08265_),
    .Y(_08287_));
 sky130_fd_sc_hd__nor2_1 _15674_ (.A(_07379_),
    .B(_08060_),
    .Y(_08288_));
 sky130_fd_sc_hd__and2b_1 _15675_ (.A_N(_08234_),
    .B(_08288_),
    .X(_08289_));
 sky130_fd_sc_hd__xnor2_1 _15676_ (.A(_08280_),
    .B(_08289_),
    .Y(_08290_));
 sky130_fd_sc_hd__xnor2_1 _15677_ (.A(_08251_),
    .B(_08260_),
    .Y(_08291_));
 sky130_fd_sc_hd__xnor2_1 _15678_ (.A(_08255_),
    .B(_08257_),
    .Y(_08292_));
 sky130_fd_sc_hd__nor2_1 _15679_ (.A(_07466_),
    .B(_07675_),
    .Y(_08293_));
 sky130_fd_sc_hd__a2bb2o_1 _15680_ (.A1_N(_07507_),
    .A2_N(_07645_),
    .B1(_08293_),
    .B2(_07882_),
    .X(_08294_));
 sky130_fd_sc_hd__and2_1 _15681_ (.A(_07481_),
    .B(_07482_),
    .X(_08295_));
 sky130_fd_sc_hd__buf_4 _15682_ (.A(_08295_),
    .X(_08296_));
 sky130_fd_sc_hd__nor2_1 _15683_ (.A(_08296_),
    .B(_07842_),
    .Y(_08297_));
 sky130_fd_sc_hd__or4_1 _15684_ (.A(_07507_),
    .B(_07879_),
    .C(_07645_),
    .D(_07718_),
    .X(_08298_));
 sky130_fd_sc_hd__a21bo_1 _15685_ (.A1(_08294_),
    .A2(_08297_),
    .B1_N(_08298_),
    .X(_08299_));
 sky130_fd_sc_hd__xnor2_1 _15686_ (.A(_08292_),
    .B(_08299_),
    .Y(_08300_));
 sky130_fd_sc_hd__nor2_1 _15687_ (.A(_08274_),
    .B(_07971_),
    .Y(_08301_));
 sky130_fd_sc_hd__xnor2_1 _15688_ (.A(_08275_),
    .B(_08301_),
    .Y(_08302_));
 sky130_fd_sc_hd__xnor2_1 _15689_ (.A(_08273_),
    .B(_08302_),
    .Y(_08303_));
 sky130_fd_sc_hd__and2b_1 _15690_ (.A_N(_08292_),
    .B(_08299_),
    .X(_08304_));
 sky130_fd_sc_hd__a21o_1 _15691_ (.A1(_08300_),
    .A2(_08303_),
    .B1(_08304_),
    .X(_08305_));
 sky130_fd_sc_hd__xnor2_1 _15692_ (.A(_08291_),
    .B(_08305_),
    .Y(_08306_));
 sky130_fd_sc_hd__or2b_1 _15693_ (.A(_08291_),
    .B_N(_08305_),
    .X(_08307_));
 sky130_fd_sc_hd__a21boi_1 _15694_ (.A1(_08290_),
    .A2(_08306_),
    .B1_N(_08307_),
    .Y(_08308_));
 sky130_fd_sc_hd__xor2_1 _15695_ (.A(_08287_),
    .B(_08308_),
    .X(_08309_));
 sky130_fd_sc_hd__nor2_1 _15696_ (.A(_08287_),
    .B(_08308_),
    .Y(_08310_));
 sky130_fd_sc_hd__a21oi_1 _15697_ (.A1(_08286_),
    .A2(_08309_),
    .B1(_08310_),
    .Y(_08311_));
 sky130_fd_sc_hd__xor2_1 _15698_ (.A(_08284_),
    .B(_08311_),
    .X(_08312_));
 sky130_fd_sc_hd__nor2_1 _15699_ (.A(_08284_),
    .B(_08311_),
    .Y(_08313_));
 sky130_fd_sc_hd__a21oi_1 _15700_ (.A1(_08283_),
    .A2(_08312_),
    .B1(_08313_),
    .Y(_08314_));
 sky130_fd_sc_hd__xnor2_2 _15701_ (.A(_08188_),
    .B(_08215_),
    .Y(_08315_));
 sky130_fd_sc_hd__nor2_1 _15702_ (.A(_08245_),
    .B(_08269_),
    .Y(_08316_));
 sky130_fd_sc_hd__a21oi_2 _15703_ (.A1(_08244_),
    .A2(_08270_),
    .B1(_08316_),
    .Y(_08317_));
 sky130_fd_sc_hd__xnor2_2 _15704_ (.A(_08315_),
    .B(_08317_),
    .Y(_08318_));
 sky130_fd_sc_hd__nor3_1 _15705_ (.A(_08271_),
    .B(_08314_),
    .C(_08318_),
    .Y(_08319_));
 sky130_fd_sc_hd__nor2_1 _15706_ (.A(_08315_),
    .B(_08317_),
    .Y(_08320_));
 sky130_fd_sc_hd__nor2_1 _15707_ (.A(_08320_),
    .B(_08319_),
    .Y(_08321_));
 sky130_fd_sc_hd__xnor2_2 _15708_ (.A(_08221_),
    .B(_08321_),
    .Y(_08322_));
 sky130_fd_sc_hd__xnor2_1 _15709_ (.A(_08286_),
    .B(_08309_),
    .Y(_08323_));
 sky130_fd_sc_hd__or4_2 _15710_ (.A(_07435_),
    .B(_08256_),
    .C(_07592_),
    .D(_07970_),
    .X(_08324_));
 sky130_fd_sc_hd__or2_1 _15711_ (.A(_07467_),
    .B(_07986_),
    .X(_08325_));
 sky130_fd_sc_hd__o22ai_1 _15712_ (.A1(_07470_),
    .A2(_07593_),
    .B1(_07971_),
    .B2(_08256_),
    .Y(_08326_));
 sky130_fd_sc_hd__and2_1 _15713_ (.A(_08324_),
    .B(_08326_),
    .X(_08327_));
 sky130_fd_sc_hd__or2b_1 _15714_ (.A(_08325_),
    .B_N(_08327_),
    .X(_08328_));
 sky130_fd_sc_hd__o22a_1 _15715_ (.A1(_08272_),
    .A2(_07986_),
    .B1(_08060_),
    .B2(_07400_),
    .X(_08329_));
 sky130_fd_sc_hd__a211oi_2 _15716_ (.A1(_08324_),
    .A2(_08328_),
    .B1(_08329_),
    .C1(_08289_),
    .Y(_08330_));
 sky130_fd_sc_hd__xnor2_1 _15717_ (.A(_08290_),
    .B(_08306_),
    .Y(_08331_));
 sky130_fd_sc_hd__xnor2_1 _15718_ (.A(_08300_),
    .B(_08303_),
    .Y(_08332_));
 sky130_fd_sc_hd__nand3_1 _15719_ (.A(_08298_),
    .B(_08294_),
    .C(_08297_),
    .Y(_08333_));
 sky130_fd_sc_hd__a21o_1 _15720_ (.A1(_08298_),
    .A2(_08294_),
    .B1(_08297_),
    .X(_08334_));
 sky130_fd_sc_hd__buf_4 _15721_ (.A(_07718_),
    .X(_08335_));
 sky130_fd_sc_hd__o22a_1 _15722_ (.A1(_07593_),
    .A2(_07646_),
    .B1(_08335_),
    .B2(_07789_),
    .X(_08336_));
 sky130_fd_sc_hd__or4_1 _15723_ (.A(_07789_),
    .B(_07593_),
    .C(_07646_),
    .D(_07718_),
    .X(_08337_));
 sky130_fd_sc_hd__o31ai_1 _15724_ (.A1(_07879_),
    .A2(_07843_),
    .A3(_08336_),
    .B1(_08337_),
    .Y(_08338_));
 sky130_fd_sc_hd__a21o_1 _15725_ (.A1(_08333_),
    .A2(_08334_),
    .B1(_08338_),
    .X(_08339_));
 sky130_fd_sc_hd__xnor2_1 _15726_ (.A(_08325_),
    .B(_08327_),
    .Y(_08340_));
 sky130_fd_sc_hd__nand3_1 _15727_ (.A(_08333_),
    .B(_08334_),
    .C(_08338_),
    .Y(_08341_));
 sky130_fd_sc_hd__a21bo_1 _15728_ (.A1(_08339_),
    .A2(_08340_),
    .B1_N(_08341_),
    .X(_08342_));
 sky130_fd_sc_hd__xnor2_1 _15729_ (.A(_08332_),
    .B(_08342_),
    .Y(_08343_));
 sky130_fd_sc_hd__o211a_1 _15730_ (.A1(_08289_),
    .A2(_08329_),
    .B1(_08328_),
    .C1(_08324_),
    .X(_08344_));
 sky130_fd_sc_hd__nor2_1 _15731_ (.A(_08330_),
    .B(_08344_),
    .Y(_08345_));
 sky130_fd_sc_hd__and2b_1 _15732_ (.A_N(_08332_),
    .B(_08342_),
    .X(_08346_));
 sky130_fd_sc_hd__a21o_1 _15733_ (.A1(_08343_),
    .A2(_08345_),
    .B1(_08346_),
    .X(_08347_));
 sky130_fd_sc_hd__xnor2_1 _15734_ (.A(_08331_),
    .B(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__and2b_1 _15735_ (.A_N(_08331_),
    .B(_08347_),
    .X(_08349_));
 sky130_fd_sc_hd__a21oi_1 _15736_ (.A1(_08330_),
    .A2(_08348_),
    .B1(_08349_),
    .Y(_08350_));
 sky130_fd_sc_hd__or2_1 _15737_ (.A(_08323_),
    .B(_08350_),
    .X(_08351_));
 sky130_fd_sc_hd__xnor2_1 _15738_ (.A(_08283_),
    .B(_08312_),
    .Y(_08352_));
 sky130_fd_sc_hd__nor2_1 _15739_ (.A(_08351_),
    .B(_08352_),
    .Y(_08353_));
 sky130_fd_sc_hd__xor2_1 _15740_ (.A(_08271_),
    .B(_08314_),
    .X(_08354_));
 sky130_fd_sc_hd__nand2_1 _15741_ (.A(_08353_),
    .B(_08354_),
    .Y(_08355_));
 sky130_fd_sc_hd__xor2_1 _15742_ (.A(_08330_),
    .B(_08348_),
    .X(_08356_));
 sky130_fd_sc_hd__xnor2_1 _15743_ (.A(_08343_),
    .B(_08345_),
    .Y(_08357_));
 sky130_fd_sc_hd__nand3_1 _15744_ (.A(_08341_),
    .B(_08339_),
    .C(_08340_),
    .Y(_08358_));
 sky130_fd_sc_hd__a21o_1 _15745_ (.A1(_08341_),
    .A2(_08339_),
    .B1(_08340_),
    .X(_08359_));
 sky130_fd_sc_hd__nor2_1 _15746_ (.A(_07468_),
    .B(_08060_),
    .Y(_08360_));
 sky130_fd_sc_hd__or4_1 _15747_ (.A(_07435_),
    .B(_08296_),
    .C(_07971_),
    .D(_07986_),
    .X(_08361_));
 sky130_fd_sc_hd__o22ai_1 _15748_ (.A1(_08296_),
    .A2(_07971_),
    .B1(_07986_),
    .B2(_07470_),
    .Y(_08362_));
 sky130_fd_sc_hd__and2_1 _15749_ (.A(_08361_),
    .B(_08362_),
    .X(_08363_));
 sky130_fd_sc_hd__xor2_1 _15750_ (.A(_08360_),
    .B(_08363_),
    .X(_08364_));
 sky130_fd_sc_hd__and4bb_1 _15751_ (.A_N(_07880_),
    .B_N(_08336_),
    .C(_08136_),
    .D(_08337_),
    .X(_08365_));
 sky130_fd_sc_hd__and4bb_1 _15752_ (.A_N(_07789_),
    .B_N(_07593_),
    .C(_07838_),
    .D(_08293_),
    .X(_08366_));
 sky130_fd_sc_hd__o22a_1 _15753_ (.A1(_07880_),
    .A2(_07843_),
    .B1(_08366_),
    .B2(_08336_),
    .X(_08367_));
 sky130_fd_sc_hd__a21o_1 _15754_ (.A1(_07529_),
    .A2(_07984_),
    .B1(_07646_),
    .X(_08368_));
 sky130_fd_sc_hd__o21a_1 _15755_ (.A1(_07517_),
    .A2(_08335_),
    .B1(_08368_),
    .X(_08369_));
 sky130_fd_sc_hd__or3_1 _15756_ (.A(_07517_),
    .B(_08335_),
    .C(_08368_),
    .X(_08370_));
 sky130_fd_sc_hd__o31a_1 _15757_ (.A1(_07792_),
    .A2(_07843_),
    .A3(_08369_),
    .B1(_08370_),
    .X(_08371_));
 sky130_fd_sc_hd__o21ai_1 _15758_ (.A1(_08365_),
    .A2(_08367_),
    .B1(_08371_),
    .Y(_08372_));
 sky130_fd_sc_hd__nor3_1 _15759_ (.A(_08365_),
    .B(_08367_),
    .C(_08371_),
    .Y(_08373_));
 sky130_fd_sc_hd__a21o_1 _15760_ (.A1(_08364_),
    .A2(_08372_),
    .B1(_08373_),
    .X(_08374_));
 sky130_fd_sc_hd__a21o_1 _15761_ (.A1(_08358_),
    .A2(_08359_),
    .B1(_08374_),
    .X(_08375_));
 sky130_fd_sc_hd__a21boi_1 _15762_ (.A1(_08360_),
    .A2(_08362_),
    .B1_N(_08361_),
    .Y(_08376_));
 sky130_fd_sc_hd__and2b_1 _15763_ (.A_N(_08376_),
    .B(_08288_),
    .X(_08377_));
 sky130_fd_sc_hd__and2b_1 _15764_ (.A_N(_08288_),
    .B(_08376_),
    .X(_08378_));
 sky130_fd_sc_hd__nor2_1 _15765_ (.A(_08377_),
    .B(_08378_),
    .Y(_08379_));
 sky130_fd_sc_hd__nand3_1 _15766_ (.A(_08358_),
    .B(_08359_),
    .C(_08374_),
    .Y(_08380_));
 sky130_fd_sc_hd__a21boi_1 _15767_ (.A1(_08375_),
    .A2(_08379_),
    .B1_N(_08380_),
    .Y(_08381_));
 sky130_fd_sc_hd__nor2_1 _15768_ (.A(_08357_),
    .B(_08381_),
    .Y(_08382_));
 sky130_fd_sc_hd__nor2_1 _15769_ (.A(_08356_),
    .B(_08382_),
    .Y(_08383_));
 sky130_fd_sc_hd__and2_1 _15770_ (.A(_08357_),
    .B(_08381_),
    .X(_08384_));
 sky130_fd_sc_hd__nor2_1 _15771_ (.A(_08382_),
    .B(_08384_),
    .Y(_08385_));
 sky130_fd_sc_hd__xnor2_1 _15772_ (.A(_08377_),
    .B(_08385_),
    .Y(_08386_));
 sky130_fd_sc_hd__and2b_1 _15773_ (.A_N(_08373_),
    .B(_08372_),
    .X(_08387_));
 sky130_fd_sc_hd__xnor2_1 _15774_ (.A(_08364_),
    .B(_08387_),
    .Y(_08388_));
 sky130_fd_sc_hd__nor2_1 _15775_ (.A(_07517_),
    .B(_08335_),
    .Y(_08389_));
 sky130_fd_sc_hd__xnor2_1 _15776_ (.A(_08368_),
    .B(_08389_),
    .Y(_08390_));
 sky130_fd_sc_hd__nor2_1 _15777_ (.A(_07792_),
    .B(_07843_),
    .Y(_08391_));
 sky130_fd_sc_hd__xnor2_1 _15778_ (.A(_08390_),
    .B(_08391_),
    .Y(_08392_));
 sky130_fd_sc_hd__nor2_1 _15779_ (.A(_07616_),
    .B(_07675_),
    .Y(_08393_));
 sky130_fd_sc_hd__o21ba_1 _15780_ (.A1(_07646_),
    .A2(_08059_),
    .B1_N(_08393_),
    .X(_08394_));
 sky130_fd_sc_hd__or3b_1 _15781_ (.A(_07645_),
    .B(_08059_),
    .C_N(_08393_),
    .X(_08395_));
 sky130_fd_sc_hd__o31a_1 _15782_ (.A1(_07788_),
    .A2(_07843_),
    .A3(_08394_),
    .B1(_08395_),
    .X(_08396_));
 sky130_fd_sc_hd__xor2_1 _15783_ (.A(_08392_),
    .B(_08396_),
    .X(_08397_));
 sky130_fd_sc_hd__clkbuf_4 _15784_ (.A(_07971_),
    .X(_08398_));
 sky130_fd_sc_hd__or4_1 _15785_ (.A(_07826_),
    .B(_07880_),
    .C(_08398_),
    .D(_08060_),
    .X(_08399_));
 sky130_fd_sc_hd__o22ai_1 _15786_ (.A1(_07880_),
    .A2(_08398_),
    .B1(_08060_),
    .B2(_07826_),
    .Y(_08400_));
 sky130_fd_sc_hd__and2_1 _15787_ (.A(_08399_),
    .B(_08400_),
    .X(_08401_));
 sky130_fd_sc_hd__nor2_1 _15788_ (.A(_08392_),
    .B(_08396_),
    .Y(_08402_));
 sky130_fd_sc_hd__a21oi_1 _15789_ (.A1(_08397_),
    .A2(_08401_),
    .B1(_08402_),
    .Y(_08403_));
 sky130_fd_sc_hd__nor2_1 _15790_ (.A(_08388_),
    .B(_08403_),
    .Y(_08404_));
 sky130_fd_sc_hd__xnor2_1 _15791_ (.A(_08388_),
    .B(_08403_),
    .Y(_08405_));
 sky130_fd_sc_hd__nor2_1 _15792_ (.A(_08399_),
    .B(_08405_),
    .Y(_08406_));
 sky130_fd_sc_hd__and3_1 _15793_ (.A(_08380_),
    .B(_08375_),
    .C(_08379_),
    .X(_08407_));
 sky130_fd_sc_hd__a21oi_1 _15794_ (.A1(_08380_),
    .A2(_08375_),
    .B1(_08379_),
    .Y(_08408_));
 sky130_fd_sc_hd__nor2_1 _15795_ (.A(_08407_),
    .B(_08408_),
    .Y(_08409_));
 sky130_fd_sc_hd__o21ai_1 _15796_ (.A1(_08404_),
    .A2(_08406_),
    .B1(_08409_),
    .Y(_08410_));
 sky130_fd_sc_hd__nor3_1 _15797_ (.A(_08383_),
    .B(_08386_),
    .C(_08410_),
    .Y(_08411_));
 sky130_fd_sc_hd__nand2_1 _15798_ (.A(_08323_),
    .B(_08350_),
    .Y(_08412_));
 sky130_fd_sc_hd__nand2_1 _15799_ (.A(_08351_),
    .B(_08412_),
    .Y(_08413_));
 sky130_fd_sc_hd__a21o_1 _15800_ (.A1(_08377_),
    .A2(_08385_),
    .B1(_08382_),
    .X(_08414_));
 sky130_fd_sc_hd__nand2_1 _15801_ (.A(_08356_),
    .B(_08414_),
    .Y(_08415_));
 sky130_fd_sc_hd__nor2_1 _15802_ (.A(_08413_),
    .B(_08415_),
    .Y(_08416_));
 sky130_fd_sc_hd__and2_1 _15803_ (.A(_08356_),
    .B(_08382_),
    .X(_08417_));
 sky130_fd_sc_hd__xnor2_1 _15804_ (.A(_08397_),
    .B(_08401_),
    .Y(_08418_));
 sky130_fd_sc_hd__or4b_1 _15805_ (.A(_07517_),
    .B(_08394_),
    .C(_07842_),
    .D_N(_08395_),
    .X(_08419_));
 sky130_fd_sc_hd__o21bai_1 _15806_ (.A1(_07835_),
    .A2(_08059_),
    .B1_N(_08393_),
    .Y(_08420_));
 sky130_fd_sc_hd__a22o_1 _15807_ (.A1(_07521_),
    .A2(_08136_),
    .B1(_08395_),
    .B2(_08420_),
    .X(_08421_));
 sky130_fd_sc_hd__and2_1 _15808_ (.A(_08419_),
    .B(_08421_),
    .X(_08422_));
 sky130_fd_sc_hd__nor4_2 _15809_ (.A(_07616_),
    .B(_07625_),
    .C(_07680_),
    .D(_07847_),
    .Y(_08423_));
 sky130_fd_sc_hd__nand2_1 _15810_ (.A(_08422_),
    .B(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__xnor2_1 _15811_ (.A(_08422_),
    .B(_08423_),
    .Y(_08425_));
 sky130_fd_sc_hd__or3_1 _15812_ (.A(_07878_),
    .B(_08398_),
    .C(_08425_),
    .X(_08426_));
 sky130_fd_sc_hd__a21o_1 _15813_ (.A1(_08424_),
    .A2(_08426_),
    .B1(_08418_),
    .X(_08427_));
 sky130_fd_sc_hd__o21a_1 _15814_ (.A1(_07878_),
    .A2(_08398_),
    .B1(_08425_),
    .X(_08428_));
 sky130_fd_sc_hd__clkbuf_4 _15815_ (.A(_07616_),
    .X(_08429_));
 sky130_fd_sc_hd__o22a_1 _15816_ (.A1(_07625_),
    .A2(_07680_),
    .B1(_07847_),
    .B2(_08429_),
    .X(_08430_));
 sky130_fd_sc_hd__a21oi_1 _15817_ (.A1(_07788_),
    .A2(_07680_),
    .B1(_08389_),
    .Y(_08431_));
 sky130_fd_sc_hd__or4_1 _15818_ (.A(_07616_),
    .B(_07633_),
    .C(_07847_),
    .D(_08431_),
    .X(_08432_));
 sky130_fd_sc_hd__o31ai_1 _15819_ (.A1(_07788_),
    .A2(_08423_),
    .A3(_08430_),
    .B1(_08432_),
    .Y(_08433_));
 sky130_fd_sc_hd__or4bb_1 _15820_ (.A(_08428_),
    .B(_08398_),
    .C_N(_08426_),
    .D_N(_08433_),
    .X(_08434_));
 sky130_fd_sc_hd__a221o_1 _15821_ (.A1(_08418_),
    .A2(_08424_),
    .B1(_08427_),
    .B2(_08434_),
    .C1(_08406_),
    .X(_08435_));
 sky130_fd_sc_hd__nand2_1 _15822_ (.A(_08399_),
    .B(_08405_),
    .Y(_08436_));
 sky130_fd_sc_hd__or2_1 _15823_ (.A(_08409_),
    .B(_08404_),
    .X(_08437_));
 sky130_fd_sc_hd__and4b_1 _15824_ (.A_N(_08435_),
    .B(_08436_),
    .C(_08410_),
    .D(_08437_),
    .X(_08438_));
 sky130_fd_sc_hd__or4b_1 _15825_ (.A(_08383_),
    .B(_08417_),
    .C(_08386_),
    .D_N(_08438_),
    .X(_08439_));
 sky130_fd_sc_hd__o21a_1 _15826_ (.A1(_08413_),
    .A2(_08439_),
    .B1(_08415_),
    .X(_08440_));
 sky130_fd_sc_hd__a21oi_1 _15827_ (.A1(_08352_),
    .A2(_08416_),
    .B1(_08440_),
    .Y(_08441_));
 sky130_fd_sc_hd__nand2_1 _15828_ (.A(_08413_),
    .B(_08439_),
    .Y(_08442_));
 sky130_fd_sc_hd__xor2_1 _15829_ (.A(_08351_),
    .B(_08352_),
    .X(_08443_));
 sky130_fd_sc_hd__o22a_1 _15830_ (.A1(_08353_),
    .A2(_08354_),
    .B1(_08416_),
    .B2(_08443_),
    .X(_08444_));
 sky130_fd_sc_hd__o2111a_1 _15831_ (.A1(_08411_),
    .A2(_08441_),
    .B1(_08355_),
    .C1(_08442_),
    .D1(_08444_),
    .X(_08445_));
 sky130_fd_sc_hd__nor2_1 _15832_ (.A(_08271_),
    .B(_08314_),
    .Y(_08446_));
 sky130_fd_sc_hd__a21o_1 _15833_ (.A1(_08353_),
    .A2(_08354_),
    .B1(_08446_),
    .X(_08447_));
 sky130_fd_sc_hd__xnor2_1 _15834_ (.A(_08318_),
    .B(_08447_),
    .Y(_08448_));
 sky130_fd_sc_hd__a2bb2o_2 _15835_ (.A1_N(_08355_),
    .A2_N(_08318_),
    .B1(_08445_),
    .B2(_08448_),
    .X(_08449_));
 sky130_fd_sc_hd__a22o_1 _15836_ (.A1(_08221_),
    .A2(_08319_),
    .B1(_08322_),
    .B2(_08449_),
    .X(_08450_));
 sky130_fd_sc_hd__xnor2_1 _15837_ (.A(_08172_),
    .B(_08218_),
    .Y(_08451_));
 sky130_fd_sc_hd__a21o_1 _15838_ (.A1(_08221_),
    .A2(_08320_),
    .B1(_08451_),
    .X(_08452_));
 sky130_fd_sc_hd__and3b_1 _15839_ (.A_N(_08172_),
    .B(_08221_),
    .C(_08320_),
    .X(_08453_));
 sky130_fd_sc_hd__a21o_1 _15840_ (.A1(_08450_),
    .A2(_08452_),
    .B1(_08453_),
    .X(_08454_));
 sky130_fd_sc_hd__nor2_1 _15841_ (.A(_08167_),
    .B(_08219_),
    .Y(_08455_));
 sky130_fd_sc_hd__xnor2_1 _15842_ (.A(_08112_),
    .B(_08455_),
    .Y(_08456_));
 sky130_fd_sc_hd__a22o_2 _15843_ (.A1(_08112_),
    .A2(_08219_),
    .B1(_08454_),
    .B2(_08456_),
    .X(_08457_));
 sky130_fd_sc_hd__a21oi_1 _15844_ (.A1(_08109_),
    .A2(_08169_),
    .B1(_08035_),
    .Y(_08458_));
 sky130_fd_sc_hd__a31o_2 _15845_ (.A1(_08110_),
    .A2(_08171_),
    .A3(_08457_),
    .B1(_08458_),
    .X(_08459_));
 sky130_fd_sc_hd__nor2_1 _15846_ (.A(_07961_),
    .B(_08034_),
    .Y(_08460_));
 sky130_fd_sc_hd__a2bb2o_1 _15847_ (.A1_N(_07863_),
    .A2_N(_07865_),
    .B1(_07748_),
    .B2(_07862_),
    .X(_08461_));
 sky130_fd_sc_hd__a21boi_1 _15848_ (.A1(_07815_),
    .A2(_07828_),
    .B1_N(_07825_),
    .Y(_08462_));
 sky130_fd_sc_hd__a21oi_1 _15849_ (.A1(_07672_),
    .A2(_07673_),
    .B1(_07379_),
    .Y(_08463_));
 sky130_fd_sc_hd__a2111o_1 _15850_ (.A1(_07672_),
    .A2(_07673_),
    .B1(_07711_),
    .C1(_07400_),
    .D1(_07379_),
    .X(_08464_));
 sky130_fd_sc_hd__o21ai_1 _15851_ (.A1(_07862_),
    .A2(_08463_),
    .B1(_08464_),
    .Y(_08465_));
 sky130_fd_sc_hd__nor2_1 _15852_ (.A(_07751_),
    .B(_07736_),
    .Y(_08466_));
 sky130_fd_sc_hd__xnor2_1 _15853_ (.A(_08465_),
    .B(_08466_),
    .Y(_08467_));
 sky130_fd_sc_hd__and2b_1 _15854_ (.A_N(_08462_),
    .B(_08467_),
    .X(_08468_));
 sky130_fd_sc_hd__and2b_1 _15855_ (.A_N(_08467_),
    .B(_08462_),
    .X(_08469_));
 sky130_fd_sc_hd__nor2_1 _15856_ (.A(_08468_),
    .B(_08469_),
    .Y(_08470_));
 sky130_fd_sc_hd__xor2_1 _15857_ (.A(_08461_),
    .B(_08470_),
    .X(_08471_));
 sky130_fd_sc_hd__nor2_1 _15858_ (.A(_07814_),
    .B(_07817_),
    .Y(_08472_));
 sky130_fd_sc_hd__nand2_1 _15859_ (.A(_07453_),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .Y(_08473_));
 sky130_fd_sc_hd__or4_2 _15860_ (.A(_07217_),
    .B(_07221_),
    .C(_07225_),
    .D(_07687_),
    .X(_08474_));
 sky130_fd_sc_hd__o211a_1 _15861_ (.A1(_07223_),
    .A2(_07096_),
    .B1(_07101_),
    .C1(_07224_),
    .X(_08475_));
 sky130_fd_sc_hd__a31o_1 _15862_ (.A1(_07689_),
    .A2(_07819_),
    .A3(_07690_),
    .B1(_08475_),
    .X(_08476_));
 sky130_fd_sc_hd__a31o_1 _15863_ (.A1(_04933_),
    .A2(_08474_),
    .A3(_08476_),
    .B1(_07822_),
    .X(_08477_));
 sky130_fd_sc_hd__a21o_2 _15864_ (.A1(_08473_),
    .A2(_08477_),
    .B1(_04937_),
    .X(_08478_));
 sky130_fd_sc_hd__or4_1 _15865_ (.A(_07470_),
    .B(_07471_),
    .C(_07834_),
    .D(_08478_),
    .X(_08479_));
 sky130_fd_sc_hd__a2bb2o_1 _15866_ (.A1_N(_07471_),
    .A2_N(_08478_),
    .B1(_07837_),
    .B2(_07697_),
    .X(_08480_));
 sky130_fd_sc_hd__and3_1 _15867_ (.A(_08472_),
    .B(_08479_),
    .C(_08480_),
    .X(_08481_));
 sky130_fd_sc_hd__a21oi_1 _15868_ (.A1(_08479_),
    .A2(_08480_),
    .B1(_08472_),
    .Y(_08482_));
 sky130_fd_sc_hd__nor2_1 _15869_ (.A(_08481_),
    .B(_08482_),
    .Y(_08483_));
 sky130_fd_sc_hd__nand2_1 _15870_ (.A(_07466_),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .Y(_08484_));
 sky130_fd_sc_hd__a21bo_1 _15871_ (.A1(_07661_),
    .A2(_07662_),
    .B1_N(_08484_),
    .X(_08485_));
 sky130_fd_sc_hd__or4b_1 _15872_ (.A(_07646_),
    .B(_07840_),
    .C(_08335_),
    .D_N(_08485_),
    .X(_08486_));
 sky130_fd_sc_hd__a2bb2o_1 _15873_ (.A1_N(_07840_),
    .A2_N(_08335_),
    .B1(_08485_),
    .B2(_07838_),
    .X(_08487_));
 sky130_fd_sc_hd__or4bb_1 _15874_ (.A(_07824_),
    .B(_07847_),
    .C_N(_08486_),
    .D_N(_08487_),
    .X(_08488_));
 sky130_fd_sc_hd__a2bb2o_1 _15875_ (.A1_N(_07827_),
    .A2_N(_07847_),
    .B1(_08486_),
    .B2(_08487_),
    .X(_08489_));
 sky130_fd_sc_hd__a21bo_1 _15876_ (.A1(_07839_),
    .A2(_07844_),
    .B1_N(_07836_),
    .X(_08490_));
 sky130_fd_sc_hd__nand3_1 _15877_ (.A(_08488_),
    .B(_08489_),
    .C(_08490_),
    .Y(_08491_));
 sky130_fd_sc_hd__a21o_1 _15878_ (.A1(_08488_),
    .A2(_08489_),
    .B1(_08490_),
    .X(_08492_));
 sky130_fd_sc_hd__nand3_1 _15879_ (.A(_08483_),
    .B(_08491_),
    .C(_08492_),
    .Y(_08493_));
 sky130_fd_sc_hd__a21o_1 _15880_ (.A1(_08491_),
    .A2(_08492_),
    .B1(_08483_),
    .X(_08494_));
 sky130_fd_sc_hd__a21bo_1 _15881_ (.A1(_07830_),
    .A2(_07851_),
    .B1_N(_07850_),
    .X(_08495_));
 sky130_fd_sc_hd__nand3_1 _15882_ (.A(_08493_),
    .B(_08494_),
    .C(_08495_),
    .Y(_08496_));
 sky130_fd_sc_hd__a21o_1 _15883_ (.A1(_08493_),
    .A2(_08494_),
    .B1(_08495_),
    .X(_08497_));
 sky130_fd_sc_hd__nand3_1 _15884_ (.A(_08471_),
    .B(_08496_),
    .C(_08497_),
    .Y(_08498_));
 sky130_fd_sc_hd__a21o_1 _15885_ (.A1(_08496_),
    .A2(_08497_),
    .B1(_08471_),
    .X(_08499_));
 sky130_fd_sc_hd__a21bo_1 _15886_ (.A1(_07857_),
    .A2(_07868_),
    .B1_N(_07856_),
    .X(_08500_));
 sky130_fd_sc_hd__nand3_1 _15887_ (.A(_08498_),
    .B(_08499_),
    .C(_08500_),
    .Y(_08501_));
 sky130_fd_sc_hd__a21o_1 _15888_ (.A1(_08498_),
    .A2(_08499_),
    .B1(_08500_),
    .X(_08502_));
 sky130_fd_sc_hd__a21o_1 _15889_ (.A1(_07888_),
    .A2(_07897_),
    .B1(_07896_),
    .X(_08503_));
 sky130_fd_sc_hd__or2b_1 _15890_ (.A(_07861_),
    .B_N(_07866_),
    .X(_08504_));
 sky130_fd_sc_hd__a21bo_1 _15891_ (.A1(_07859_),
    .A2(_07867_),
    .B1_N(_08504_),
    .X(_08505_));
 sky130_fd_sc_hd__or4_1 _15892_ (.A(_07424_),
    .B(_08296_),
    .C(_07591_),
    .D(_07790_),
    .X(_08506_));
 sky130_fd_sc_hd__clkinv_2 _15893_ (.A(_08296_),
    .Y(_08507_));
 sky130_fd_sc_hd__a2bb2o_1 _15894_ (.A1_N(_07424_),
    .A2_N(_08067_),
    .B1(_07520_),
    .B2(_08507_),
    .X(_08508_));
 sky130_fd_sc_hd__nand2_1 _15895_ (.A(_08506_),
    .B(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__clkbuf_4 _15896_ (.A(_07880_),
    .X(_08510_));
 sky130_fd_sc_hd__nor2_1 _15897_ (.A(_07598_),
    .B(_08510_),
    .Y(_08511_));
 sky130_fd_sc_hd__xnor2_2 _15898_ (.A(_08509_),
    .B(_08511_),
    .Y(_08512_));
 sky130_fd_sc_hd__or4_1 _15899_ (.A(_07442_),
    .B(_07355_),
    .C(_07552_),
    .D(_07550_),
    .X(_08513_));
 sky130_fd_sc_hd__o22ai_1 _15900_ (.A1(_07742_),
    .A2(_07890_),
    .B1(_07800_),
    .B2(_07469_),
    .Y(_08514_));
 sky130_fd_sc_hd__nand2_1 _15901_ (.A(_08513_),
    .B(_08514_),
    .Y(_08515_));
 sky130_fd_sc_hd__or2_1 _15902_ (.A(_07388_),
    .B(_07567_),
    .X(_08516_));
 sky130_fd_sc_hd__xnor2_1 _15903_ (.A(_08515_),
    .B(_08516_),
    .Y(_08517_));
 sky130_fd_sc_hd__o31a_1 _15904_ (.A1(_07424_),
    .A2(_07805_),
    .A3(_07892_),
    .B1(_07889_),
    .X(_08518_));
 sky130_fd_sc_hd__nor2_1 _15905_ (.A(_08517_),
    .B(_08518_),
    .Y(_08519_));
 sky130_fd_sc_hd__nand2_1 _15906_ (.A(_08517_),
    .B(_08518_),
    .Y(_08520_));
 sky130_fd_sc_hd__and2b_1 _15907_ (.A_N(_08519_),
    .B(_08520_),
    .X(_08521_));
 sky130_fd_sc_hd__xor2_2 _15908_ (.A(_08512_),
    .B(_08521_),
    .X(_08522_));
 sky130_fd_sc_hd__xnor2_1 _15909_ (.A(_08505_),
    .B(_08522_),
    .Y(_08523_));
 sky130_fd_sc_hd__xnor2_1 _15910_ (.A(_08503_),
    .B(_08523_),
    .Y(_08524_));
 sky130_fd_sc_hd__and3_1 _15911_ (.A(_08501_),
    .B(_08502_),
    .C(_08524_),
    .X(_08525_));
 sky130_fd_sc_hd__a21oi_1 _15912_ (.A1(_08501_),
    .A2(_08502_),
    .B1(_08524_),
    .Y(_08526_));
 sky130_fd_sc_hd__or2_1 _15913_ (.A(_08525_),
    .B(_08526_),
    .X(_08527_));
 sky130_fd_sc_hd__and2_1 _15914_ (.A(_07873_),
    .B(_07904_),
    .X(_08528_));
 sky130_fd_sc_hd__xor2_1 _15915_ (.A(_08527_),
    .B(_08528_),
    .X(_08529_));
 sky130_fd_sc_hd__or2b_1 _15916_ (.A(_07902_),
    .B_N(_07875_),
    .X(_08530_));
 sky130_fd_sc_hd__nand2_4 _15917_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_03796_),
    .Y(_08531_));
 sky130_fd_sc_hd__nor2_1 _15918_ (.A(_07625_),
    .B(_08531_),
    .Y(_08532_));
 sky130_fd_sc_hd__a21o_1 _15919_ (.A1(_07913_),
    .A2(_07917_),
    .B1(_07911_),
    .X(_08533_));
 sky130_fd_sc_hd__inv_2 _15920_ (.A(_08533_),
    .Y(_08534_));
 sky130_fd_sc_hd__or4b_1 _15921_ (.A(_07792_),
    .B(_07517_),
    .C(_07620_),
    .D_N(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_08535_));
 sky130_fd_sc_hd__nor2_2 _15922_ (.A(_04938_),
    .B(_07617_),
    .Y(_08536_));
 sky130_fd_sc_hd__a2bb2o_1 _15923_ (.A1_N(_07792_),
    .A2_N(_07621_),
    .B1(_08536_),
    .B2(_07521_),
    .X(_08537_));
 sky130_fd_sc_hd__nand2_1 _15924_ (.A(_08535_),
    .B(_08537_),
    .Y(_08538_));
 sky130_fd_sc_hd__nor2_1 _15925_ (.A(_07616_),
    .B(_07914_),
    .Y(_08539_));
 sky130_fd_sc_hd__xor2_1 _15926_ (.A(_08538_),
    .B(_08539_),
    .X(_08540_));
 sky130_fd_sc_hd__a21o_1 _15927_ (.A1(_07881_),
    .A2(_07885_),
    .B1(_08540_),
    .X(_08541_));
 sky130_fd_sc_hd__nand3_1 _15928_ (.A(_07881_),
    .B(_07885_),
    .C(_08540_),
    .Y(_08542_));
 sky130_fd_sc_hd__nand2_1 _15929_ (.A(_08541_),
    .B(_08542_),
    .Y(_08543_));
 sky130_fd_sc_hd__xnor2_1 _15930_ (.A(_08534_),
    .B(_08543_),
    .Y(_08544_));
 sky130_fd_sc_hd__o21bai_1 _15931_ (.A1(_07623_),
    .A2(_07920_),
    .B1_N(_07919_),
    .Y(_08545_));
 sky130_fd_sc_hd__xor2_1 _15932_ (.A(_08544_),
    .B(_08545_),
    .X(_08546_));
 sky130_fd_sc_hd__xnor2_1 _15933_ (.A(_08532_),
    .B(_08546_),
    .Y(_08547_));
 sky130_fd_sc_hd__a21o_1 _15934_ (.A1(_07900_),
    .A2(_08530_),
    .B1(_08547_),
    .X(_08548_));
 sky130_fd_sc_hd__nand3_1 _15935_ (.A(_07900_),
    .B(_08530_),
    .C(_08547_),
    .Y(_08549_));
 sky130_fd_sc_hd__nand2_1 _15936_ (.A(_08548_),
    .B(_08549_),
    .Y(_08550_));
 sky130_fd_sc_hd__nor2_1 _15937_ (.A(_07628_),
    .B(_07921_),
    .Y(_08551_));
 sky130_fd_sc_hd__xnor2_2 _15938_ (.A(_08550_),
    .B(_08551_),
    .Y(_08552_));
 sky130_fd_sc_hd__xnor2_1 _15939_ (.A(_08529_),
    .B(_08552_),
    .Y(_08553_));
 sky130_fd_sc_hd__and2_1 _15940_ (.A(_07906_),
    .B(_07928_),
    .X(_08554_));
 sky130_fd_sc_hd__xnor2_1 _15941_ (.A(_08553_),
    .B(_08554_),
    .Y(_08555_));
 sky130_fd_sc_hd__o21ba_1 _15942_ (.A1(_07637_),
    .A2(_07925_),
    .B1_N(_07924_),
    .X(_08556_));
 sky130_fd_sc_hd__xnor2_1 _15943_ (.A(_08555_),
    .B(_08556_),
    .Y(_08557_));
 sky130_fd_sc_hd__and3_1 _15944_ (.A(_07928_),
    .B(_07929_),
    .C(_07959_),
    .X(_08558_));
 sky130_fd_sc_hd__a21oi_1 _15945_ (.A1(_07640_),
    .A2(_07960_),
    .B1(_08558_),
    .Y(_08559_));
 sky130_fd_sc_hd__xor2_1 _15946_ (.A(_08557_),
    .B(_08559_),
    .X(_08560_));
 sky130_fd_sc_hd__nand2_1 _15947_ (.A(_08460_),
    .B(_08560_),
    .Y(_08561_));
 sky130_fd_sc_hd__or2_1 _15948_ (.A(_08460_),
    .B(_08560_),
    .X(_08562_));
 sky130_fd_sc_hd__and2_2 _15949_ (.A(_08561_),
    .B(_08562_),
    .X(_08563_));
 sky130_fd_sc_hd__xor2_2 _15950_ (.A(_08459_),
    .B(_08563_),
    .X(_08564_));
 sky130_fd_sc_hd__or2b_1 _15951_ (.A(_07344_),
    .B_N(_08564_),
    .X(_08565_));
 sky130_fd_sc_hd__or2b_1 _15952_ (.A(_08564_),
    .B_N(_07344_),
    .X(_08566_));
 sky130_fd_sc_hd__nand2_1 _15953_ (.A(_08565_),
    .B(_08566_),
    .Y(_08567_));
 sky130_fd_sc_hd__a21boi_2 _15954_ (.A1(_08171_),
    .A2(_08457_),
    .B1_N(_08169_),
    .Y(_08568_));
 sky130_fd_sc_hd__or2_1 _15955_ (.A(_08035_),
    .B(_08109_),
    .X(_08569_));
 sky130_fd_sc_hd__and2_1 _15956_ (.A(_08110_),
    .B(_08569_),
    .X(_08570_));
 sky130_fd_sc_hd__xnor2_4 _15957_ (.A(_08568_),
    .B(_08570_),
    .Y(_08571_));
 sky130_fd_sc_hd__mux2_1 _15958_ (.A0(\rbzero.debug_overlay.playerY[-7] ),
    .A1(\rbzero.debug_overlay.playerX[-7] ),
    .S(_07343_),
    .X(_08572_));
 sky130_fd_sc_hd__xnor2_4 _15959_ (.A(_08171_),
    .B(_08457_),
    .Y(_08573_));
 sky130_fd_sc_hd__inv_2 _15960_ (.A(\rbzero.debug_overlay.playerY[-8] ),
    .Y(_08574_));
 sky130_fd_sc_hd__mux2_1 _15961_ (.A0(_08574_),
    .A1(_07431_),
    .S(_07343_),
    .X(_08575_));
 sky130_fd_sc_hd__xor2_2 _15962_ (.A(_08454_),
    .B(_08456_),
    .X(_08576_));
 sky130_fd_sc_hd__mux2_1 _15963_ (.A0(\rbzero.debug_overlay.playerY[-9] ),
    .A1(\rbzero.debug_overlay.playerX[-9] ),
    .S(_07342_),
    .X(_08577_));
 sky130_fd_sc_hd__nand2_1 _15964_ (.A(_08576_),
    .B(_08577_),
    .Y(_08578_));
 sky130_fd_sc_hd__a21oi_1 _15965_ (.A1(_08573_),
    .A2(_08575_),
    .B1(_08578_),
    .Y(_08579_));
 sky130_fd_sc_hd__nor2_1 _15966_ (.A(_08573_),
    .B(_08575_),
    .Y(_08580_));
 sky130_fd_sc_hd__a211o_1 _15967_ (.A1(_08571_),
    .A2(_08572_),
    .B1(_08579_),
    .C1(_08580_),
    .X(_08581_));
 sky130_fd_sc_hd__o21ai_2 _15968_ (.A1(_08571_),
    .A2(_08572_),
    .B1(_08581_),
    .Y(_08582_));
 sky130_fd_sc_hd__xor2_1 _15969_ (.A(_08567_),
    .B(_08582_),
    .X(_08583_));
 sky130_fd_sc_hd__or2_1 _15970_ (.A(_07343_),
    .B(_07491_),
    .X(_08584_));
 sky130_fd_sc_hd__o21ai_4 _15971_ (.A1(_07334_),
    .A2(_05114_),
    .B1(_08584_),
    .Y(_08585_));
 sky130_fd_sc_hd__xnor2_1 _15972_ (.A(_08583_),
    .B(_08585_),
    .Y(_08586_));
 sky130_fd_sc_hd__nand2_1 _15973_ (.A(_07338_),
    .B(_08586_),
    .Y(_08587_));
 sky130_fd_sc_hd__o211a_1 _15974_ (.A1(\rbzero.wall_tracer.texu[0] ),
    .A2(_07338_),
    .B1(_07266_),
    .C1(_08587_),
    .X(_00481_));
 sky130_fd_sc_hd__a21boi_2 _15975_ (.A1(_08459_),
    .A2(_08563_),
    .B1_N(_08561_),
    .Y(_08588_));
 sky130_fd_sc_hd__or2_1 _15976_ (.A(_08557_),
    .B(_08559_),
    .X(_08589_));
 sky130_fd_sc_hd__a21o_1 _15977_ (.A1(_08512_),
    .A2(_08520_),
    .B1(_08519_),
    .X(_08590_));
 sky130_fd_sc_hd__a21o_1 _15978_ (.A1(_08461_),
    .A2(_08470_),
    .B1(_08468_),
    .X(_08591_));
 sky130_fd_sc_hd__clkbuf_2 _15979_ (.A(_08256_),
    .X(_08592_));
 sky130_fd_sc_hd__or4_1 _15980_ (.A(_07388_),
    .B(_08592_),
    .C(_08067_),
    .D(_07790_),
    .X(_08593_));
 sky130_fd_sc_hd__clkbuf_4 _15981_ (.A(_08067_),
    .X(_08594_));
 sky130_fd_sc_hd__clkbuf_4 _15982_ (.A(_07790_),
    .X(_08595_));
 sky130_fd_sc_hd__buf_2 _15983_ (.A(_08592_),
    .X(_08596_));
 sky130_fd_sc_hd__o22ai_1 _15984_ (.A1(_07388_),
    .A2(_08594_),
    .B1(_08595_),
    .B2(_08596_),
    .Y(_08597_));
 sky130_fd_sc_hd__nand2_1 _15985_ (.A(_08593_),
    .B(_08597_),
    .Y(_08598_));
 sky130_fd_sc_hd__buf_2 _15986_ (.A(_08296_),
    .X(_08599_));
 sky130_fd_sc_hd__nor2_1 _15987_ (.A(_08599_),
    .B(_07598_),
    .Y(_08600_));
 sky130_fd_sc_hd__xnor2_2 _15988_ (.A(_08598_),
    .B(_08600_),
    .Y(_08601_));
 sky130_fd_sc_hd__or4_1 _15989_ (.A(_07742_),
    .B(_07552_),
    .C(_07550_),
    .D(_07736_),
    .X(_08602_));
 sky130_fd_sc_hd__or2_1 _15990_ (.A(_07552_),
    .B(_07736_),
    .X(_08603_));
 sky130_fd_sc_hd__o21ai_1 _15991_ (.A1(_07742_),
    .A2(_07800_),
    .B1(_08603_),
    .Y(_08604_));
 sky130_fd_sc_hd__nand2_1 _15992_ (.A(_08602_),
    .B(_08604_),
    .Y(_08605_));
 sky130_fd_sc_hd__or2_1 _15993_ (.A(_07469_),
    .B(_07805_),
    .X(_08606_));
 sky130_fd_sc_hd__xnor2_1 _15994_ (.A(_08605_),
    .B(_08606_),
    .Y(_08607_));
 sky130_fd_sc_hd__o31a_1 _15995_ (.A1(_07388_),
    .A2(_07805_),
    .A3(_08515_),
    .B1(_08513_),
    .X(_08608_));
 sky130_fd_sc_hd__nor2_1 _15996_ (.A(_08607_),
    .B(_08608_),
    .Y(_08609_));
 sky130_fd_sc_hd__nand2_1 _15997_ (.A(_08607_),
    .B(_08608_),
    .Y(_08610_));
 sky130_fd_sc_hd__and2b_1 _15998_ (.A_N(_08609_),
    .B(_08610_),
    .X(_08611_));
 sky130_fd_sc_hd__xor2_2 _15999_ (.A(_08601_),
    .B(_08611_),
    .X(_08612_));
 sky130_fd_sc_hd__xnor2_1 _16000_ (.A(_08591_),
    .B(_08612_),
    .Y(_08613_));
 sky130_fd_sc_hd__xnor2_1 _16001_ (.A(_08590_),
    .B(_08613_),
    .Y(_08614_));
 sky130_fd_sc_hd__o31ai_1 _16002_ (.A1(_07858_),
    .A2(_07736_),
    .A3(_08465_),
    .B1(_08464_),
    .Y(_08615_));
 sky130_fd_sc_hd__a21bo_1 _16003_ (.A1(_08472_),
    .A2(_08480_),
    .B1_N(_08479_),
    .X(_08616_));
 sky130_fd_sc_hd__a21oi_2 _16004_ (.A1(_07472_),
    .A2(_07641_),
    .B1(_07400_),
    .Y(_08617_));
 sky130_fd_sc_hd__a21o_1 _16005_ (.A1(_07472_),
    .A2(_07641_),
    .B1(_07379_),
    .X(_08618_));
 sky130_fd_sc_hd__a21o_1 _16006_ (.A1(_07672_),
    .A2(_07673_),
    .B1(_07400_),
    .X(_08619_));
 sky130_fd_sc_hd__a22o_1 _16007_ (.A1(_08463_),
    .A2(_08617_),
    .B1(_08618_),
    .B2(_08619_),
    .X(_08620_));
 sky130_fd_sc_hd__nor2_1 _16008_ (.A(_07751_),
    .B(_07712_),
    .Y(_08621_));
 sky130_fd_sc_hd__xnor2_1 _16009_ (.A(_08620_),
    .B(_08621_),
    .Y(_08622_));
 sky130_fd_sc_hd__xor2_1 _16010_ (.A(_08616_),
    .B(_08622_),
    .X(_08623_));
 sky130_fd_sc_hd__nand2_1 _16011_ (.A(_08615_),
    .B(_08623_),
    .Y(_08624_));
 sky130_fd_sc_hd__or2_1 _16012_ (.A(_08615_),
    .B(_08623_),
    .X(_08625_));
 sky130_fd_sc_hd__and2_1 _16013_ (.A(_08624_),
    .B(_08625_),
    .X(_08626_));
 sky130_fd_sc_hd__nor2_1 _16014_ (.A(_07814_),
    .B(_07834_),
    .Y(_08627_));
 sky130_fd_sc_hd__and2_2 _16015_ (.A(_07663_),
    .B(_08484_),
    .X(_08628_));
 sky130_fd_sc_hd__clkbuf_4 _16016_ (.A(_07453_),
    .X(_08629_));
 sky130_fd_sc_hd__and4_1 _16017_ (.A(_07689_),
    .B(_07819_),
    .C(_08475_),
    .D(_07690_),
    .X(_08630_));
 sky130_fd_sc_hd__o41a_1 _16018_ (.A1(_07217_),
    .A2(_07221_),
    .A3(_07225_),
    .A4(_07687_),
    .B1(_07229_),
    .X(_08631_));
 sky130_fd_sc_hd__a211o_1 _16019_ (.A1(_07228_),
    .A2(_08630_),
    .B1(_08631_),
    .C1(_07337_),
    .X(_08632_));
 sky130_fd_sc_hd__a22o_4 _16020_ (.A1(_08629_),
    .A2(\rbzero.wall_tracer.stepDistY[7] ),
    .B1(_07694_),
    .B2(_08632_),
    .X(_08633_));
 sky130_fd_sc_hd__nand2_4 _16021_ (.A(_04929_),
    .B(_08633_),
    .Y(_08634_));
 sky130_fd_sc_hd__or4_1 _16022_ (.A(_07826_),
    .B(_07471_),
    .C(_08628_),
    .D(_08634_),
    .X(_08635_));
 sky130_fd_sc_hd__buf_2 _16023_ (.A(_08485_),
    .X(_08636_));
 sky130_fd_sc_hd__a32o_1 _16024_ (.A1(_04929_),
    .A2(_07698_),
    .A3(_08633_),
    .B1(_08636_),
    .B2(_07697_),
    .X(_08637_));
 sky130_fd_sc_hd__nand2_1 _16025_ (.A(_08635_),
    .B(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__xnor2_2 _16026_ (.A(_08627_),
    .B(_08638_),
    .Y(_08639_));
 sky130_fd_sc_hd__nand2_2 _16027_ (.A(_07519_),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .Y(_08640_));
 sky130_fd_sc_hd__a21oi_1 _16028_ (.A1(_07696_),
    .A2(_08640_),
    .B1(_07835_),
    .Y(_08641_));
 sky130_fd_sc_hd__nor2_1 _16029_ (.A(_07824_),
    .B(_07680_),
    .Y(_08642_));
 sky130_fd_sc_hd__xnor2_1 _16030_ (.A(_08641_),
    .B(_08642_),
    .Y(_08643_));
 sky130_fd_sc_hd__and2_1 _16031_ (.A(_08473_),
    .B(_08477_),
    .X(_08644_));
 sky130_fd_sc_hd__buf_4 _16032_ (.A(_08644_),
    .X(_08645_));
 sky130_fd_sc_hd__nor2_1 _16033_ (.A(_07843_),
    .B(_08645_),
    .Y(_08646_));
 sky130_fd_sc_hd__xor2_1 _16034_ (.A(_08643_),
    .B(_08646_),
    .X(_08647_));
 sky130_fd_sc_hd__and2_1 _16035_ (.A(_08486_),
    .B(_08488_),
    .X(_08648_));
 sky130_fd_sc_hd__xor2_1 _16036_ (.A(_08647_),
    .B(_08648_),
    .X(_08649_));
 sky130_fd_sc_hd__xnor2_2 _16037_ (.A(_08639_),
    .B(_08649_),
    .Y(_08650_));
 sky130_fd_sc_hd__and2_1 _16038_ (.A(_08491_),
    .B(_08493_),
    .X(_08651_));
 sky130_fd_sc_hd__xor2_1 _16039_ (.A(_08650_),
    .B(_08651_),
    .X(_08652_));
 sky130_fd_sc_hd__xnor2_1 _16040_ (.A(_08626_),
    .B(_08652_),
    .Y(_08653_));
 sky130_fd_sc_hd__and2_1 _16041_ (.A(_08496_),
    .B(_08498_),
    .X(_08654_));
 sky130_fd_sc_hd__xor2_1 _16042_ (.A(_08653_),
    .B(_08654_),
    .X(_08655_));
 sky130_fd_sc_hd__xnor2_1 _16043_ (.A(_08614_),
    .B(_08655_),
    .Y(_08656_));
 sky130_fd_sc_hd__a21boi_1 _16044_ (.A1(_08502_),
    .A2(_08524_),
    .B1_N(_08501_),
    .Y(_08657_));
 sky130_fd_sc_hd__xor2_1 _16045_ (.A(_08656_),
    .B(_08657_),
    .X(_08658_));
 sky130_fd_sc_hd__a2bb2o_1 _16046_ (.A1_N(_08544_),
    .A2_N(_08545_),
    .B1(_08546_),
    .B2(_08532_),
    .X(_08659_));
 sky130_fd_sc_hd__or2b_1 _16047_ (.A(_08523_),
    .B_N(_08503_),
    .X(_08660_));
 sky130_fd_sc_hd__a21bo_1 _16048_ (.A1(_08505_),
    .A2(_08522_),
    .B1_N(_08660_),
    .X(_08661_));
 sky130_fd_sc_hd__or2_1 _16049_ (.A(_08429_),
    .B(_08531_),
    .X(_08662_));
 sky130_fd_sc_hd__nand2_2 _16050_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_03796_),
    .Y(_08663_));
 sky130_fd_sc_hd__or3_2 _16051_ (.A(_07633_),
    .B(_08662_),
    .C(_08663_),
    .X(_08664_));
 sky130_fd_sc_hd__o21ai_1 _16052_ (.A1(_07633_),
    .A2(_08663_),
    .B1(_08662_),
    .Y(_08665_));
 sky130_fd_sc_hd__nand2_1 _16053_ (.A(_08664_),
    .B(_08665_),
    .Y(_08666_));
 sky130_fd_sc_hd__a21bo_1 _16054_ (.A1(_08537_),
    .A2(_08539_),
    .B1_N(_08535_),
    .X(_08667_));
 sky130_fd_sc_hd__or3b_1 _16055_ (.A(_07880_),
    .B(_07620_),
    .C_N(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_08668_));
 sky130_fd_sc_hd__or2_1 _16056_ (.A(_07792_),
    .B(_08668_),
    .X(_08669_));
 sky130_fd_sc_hd__or2_1 _16057_ (.A(_04937_),
    .B(_07617_),
    .X(_08670_));
 sky130_fd_sc_hd__clkbuf_4 _16058_ (.A(_08670_),
    .X(_08671_));
 sky130_fd_sc_hd__o22ai_1 _16059_ (.A1(_07880_),
    .A2(_07621_),
    .B1(_08671_),
    .B2(_07792_),
    .Y(_08672_));
 sky130_fd_sc_hd__nand2_1 _16060_ (.A(_08669_),
    .B(_08672_),
    .Y(_08673_));
 sky130_fd_sc_hd__nor2_1 _16061_ (.A(_07788_),
    .B(_07916_),
    .Y(_08674_));
 sky130_fd_sc_hd__xor2_1 _16062_ (.A(_08673_),
    .B(_08674_),
    .X(_08675_));
 sky130_fd_sc_hd__a21bo_1 _16063_ (.A1(_08508_),
    .A2(_08511_),
    .B1_N(_08506_),
    .X(_08676_));
 sky130_fd_sc_hd__and2b_1 _16064_ (.A_N(_08675_),
    .B(_08676_),
    .X(_08677_));
 sky130_fd_sc_hd__and2b_1 _16065_ (.A_N(_08676_),
    .B(_08675_),
    .X(_08678_));
 sky130_fd_sc_hd__nor2_1 _16066_ (.A(_08677_),
    .B(_08678_),
    .Y(_08679_));
 sky130_fd_sc_hd__xnor2_1 _16067_ (.A(_08667_),
    .B(_08679_),
    .Y(_08680_));
 sky130_fd_sc_hd__o21a_1 _16068_ (.A1(_08534_),
    .A2(_08543_),
    .B1(_08541_),
    .X(_08681_));
 sky130_fd_sc_hd__xor2_1 _16069_ (.A(_08680_),
    .B(_08681_),
    .X(_08682_));
 sky130_fd_sc_hd__xnor2_1 _16070_ (.A(_08666_),
    .B(_08682_),
    .Y(_08683_));
 sky130_fd_sc_hd__xnor2_1 _16071_ (.A(_08661_),
    .B(_08683_),
    .Y(_08684_));
 sky130_fd_sc_hd__xnor2_1 _16072_ (.A(_08659_),
    .B(_08684_),
    .Y(_08685_));
 sky130_fd_sc_hd__xnor2_1 _16073_ (.A(_08658_),
    .B(_08685_),
    .Y(_08686_));
 sky130_fd_sc_hd__nor2_1 _16074_ (.A(_08527_),
    .B(_08528_),
    .Y(_08687_));
 sky130_fd_sc_hd__a21oi_1 _16075_ (.A1(_08529_),
    .A2(_08552_),
    .B1(_08687_),
    .Y(_08688_));
 sky130_fd_sc_hd__or2_1 _16076_ (.A(_08686_),
    .B(_08688_),
    .X(_08689_));
 sky130_fd_sc_hd__nand2_1 _16077_ (.A(_08686_),
    .B(_08688_),
    .Y(_08690_));
 sky130_fd_sc_hd__nand2_1 _16078_ (.A(_08689_),
    .B(_08690_),
    .Y(_08691_));
 sky130_fd_sc_hd__o31a_1 _16079_ (.A1(_07628_),
    .A2(_07921_),
    .A3(_08550_),
    .B1(_08548_),
    .X(_08692_));
 sky130_fd_sc_hd__xnor2_1 _16080_ (.A(_08691_),
    .B(_08692_),
    .Y(_08693_));
 sky130_fd_sc_hd__or2_1 _16081_ (.A(_08553_),
    .B(_08554_),
    .X(_08694_));
 sky130_fd_sc_hd__o21a_1 _16082_ (.A1(_08555_),
    .A2(_08556_),
    .B1(_08694_),
    .X(_08695_));
 sky130_fd_sc_hd__xnor2_1 _16083_ (.A(_08693_),
    .B(_08695_),
    .Y(_08696_));
 sky130_fd_sc_hd__or2_1 _16084_ (.A(_08589_),
    .B(_08696_),
    .X(_08697_));
 sky130_fd_sc_hd__nand2_1 _16085_ (.A(_08589_),
    .B(_08696_),
    .Y(_08698_));
 sky130_fd_sc_hd__nand2_2 _16086_ (.A(_08697_),
    .B(_08698_),
    .Y(_08699_));
 sky130_fd_sc_hd__xnor2_4 _16087_ (.A(_08588_),
    .B(_08699_),
    .Y(_08700_));
 sky130_fd_sc_hd__mux2_1 _16088_ (.A0(_07389_),
    .A1(_07394_),
    .S(_07343_),
    .X(_08701_));
 sky130_fd_sc_hd__nor2_1 _16089_ (.A(_08700_),
    .B(_08701_),
    .Y(_08702_));
 sky130_fd_sc_hd__and2_1 _16090_ (.A(_08700_),
    .B(_08701_),
    .X(_08703_));
 sky130_fd_sc_hd__or2_1 _16091_ (.A(_08702_),
    .B(_08703_),
    .X(_08704_));
 sky130_fd_sc_hd__o21a_1 _16092_ (.A1(_08567_),
    .A2(_08582_),
    .B1(_08565_),
    .X(_08705_));
 sky130_fd_sc_hd__xnor2_1 _16093_ (.A(_08704_),
    .B(_08705_),
    .Y(_08706_));
 sky130_fd_sc_hd__nor2_1 _16094_ (.A(_08585_),
    .B(_08706_),
    .Y(_08707_));
 sky130_fd_sc_hd__a21o_1 _16095_ (.A1(_08585_),
    .A2(_08706_),
    .B1(_04933_),
    .X(_08708_));
 sky130_fd_sc_hd__o221a_1 _16096_ (.A1(\rbzero.wall_tracer.texu[1] ),
    .A2(_07338_),
    .B1(_08707_),
    .B2(_08708_),
    .C1(_07266_),
    .X(_00482_));
 sky130_fd_sc_hd__a21oi_1 _16097_ (.A1(_08589_),
    .A2(_08561_),
    .B1(_08696_),
    .Y(_08709_));
 sky130_fd_sc_hd__a41o_2 _16098_ (.A1(_08459_),
    .A2(_08563_),
    .A3(_08697_),
    .A4(_08698_),
    .B1(_08709_),
    .X(_08710_));
 sky130_fd_sc_hd__nor2_1 _16099_ (.A(_08693_),
    .B(_08695_),
    .Y(_08711_));
 sky130_fd_sc_hd__or2b_1 _16100_ (.A(_08666_),
    .B_N(_08682_),
    .X(_08712_));
 sky130_fd_sc_hd__o21ai_1 _16101_ (.A1(_08680_),
    .A2(_08681_),
    .B1(_08712_),
    .Y(_08713_));
 sky130_fd_sc_hd__or2b_1 _16102_ (.A(_08613_),
    .B_N(_08590_),
    .X(_08714_));
 sky130_fd_sc_hd__a21bo_1 _16103_ (.A1(_08591_),
    .A2(_08612_),
    .B1_N(_08714_),
    .X(_08715_));
 sky130_fd_sc_hd__or2_1 _16104_ (.A(_07519_),
    .B(_08531_),
    .X(_08716_));
 sky130_fd_sc_hd__buf_2 _16105_ (.A(_08716_),
    .X(_08717_));
 sky130_fd_sc_hd__buf_2 _16106_ (.A(_08717_),
    .X(_08718_));
 sky130_fd_sc_hd__or4_1 _16107_ (.A(_07788_),
    .B(_07616_),
    .C(_08718_),
    .D(_08663_),
    .X(_08719_));
 sky130_fd_sc_hd__o22ai_1 _16108_ (.A1(_07788_),
    .A2(_08718_),
    .B1(_08663_),
    .B2(_08429_),
    .Y(_08720_));
 sky130_fd_sc_hd__nand2_1 _16109_ (.A(_08719_),
    .B(_08720_),
    .Y(_08721_));
 sky130_fd_sc_hd__or3_1 _16110_ (.A(_05290_),
    .B(_08629_),
    .C(_04938_),
    .X(_08722_));
 sky130_fd_sc_hd__clkbuf_4 _16111_ (.A(_08722_),
    .X(_08723_));
 sky130_fd_sc_hd__clkbuf_4 _16112_ (.A(_08723_),
    .X(_08724_));
 sky130_fd_sc_hd__clkbuf_4 _16113_ (.A(_08724_),
    .X(_08725_));
 sky130_fd_sc_hd__nor2_1 _16114_ (.A(_07625_),
    .B(_08725_),
    .Y(_08726_));
 sky130_fd_sc_hd__xnor2_1 _16115_ (.A(_08721_),
    .B(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__xnor2_1 _16116_ (.A(_08664_),
    .B(_08727_),
    .Y(_08728_));
 sky130_fd_sc_hd__a21bo_1 _16117_ (.A1(_08672_),
    .A2(_08674_),
    .B1_N(_08669_),
    .X(_08729_));
 sky130_fd_sc_hd__a21bo_1 _16118_ (.A1(_08597_),
    .A2(_08600_),
    .B1_N(_08593_),
    .X(_08730_));
 sky130_fd_sc_hd__or2_1 _16119_ (.A(_08599_),
    .B(_08668_),
    .X(_08731_));
 sky130_fd_sc_hd__buf_2 _16120_ (.A(_07621_),
    .X(_08732_));
 sky130_fd_sc_hd__a2bb2o_1 _16121_ (.A1_N(_08599_),
    .A2_N(_08732_),
    .B1(_08536_),
    .B2(_07882_),
    .X(_08733_));
 sky130_fd_sc_hd__nand2_1 _16122_ (.A(_08731_),
    .B(_08733_),
    .Y(_08734_));
 sky130_fd_sc_hd__clkbuf_4 _16123_ (.A(_07916_),
    .X(_08735_));
 sky130_fd_sc_hd__nor2_1 _16124_ (.A(_07878_),
    .B(_08735_),
    .Y(_08736_));
 sky130_fd_sc_hd__xor2_1 _16125_ (.A(_08734_),
    .B(_08736_),
    .X(_08737_));
 sky130_fd_sc_hd__xnor2_1 _16126_ (.A(_08730_),
    .B(_08737_),
    .Y(_08738_));
 sky130_fd_sc_hd__xnor2_1 _16127_ (.A(_08729_),
    .B(_08738_),
    .Y(_08739_));
 sky130_fd_sc_hd__a21oi_1 _16128_ (.A1(_08667_),
    .A2(_08679_),
    .B1(_08677_),
    .Y(_08740_));
 sky130_fd_sc_hd__nor2_1 _16129_ (.A(_08739_),
    .B(_08740_),
    .Y(_08741_));
 sky130_fd_sc_hd__and2_1 _16130_ (.A(_08739_),
    .B(_08740_),
    .X(_08742_));
 sky130_fd_sc_hd__nor2_1 _16131_ (.A(_08741_),
    .B(_08742_),
    .Y(_08743_));
 sky130_fd_sc_hd__xor2_1 _16132_ (.A(_08728_),
    .B(_08743_),
    .X(_08744_));
 sky130_fd_sc_hd__xnor2_1 _16133_ (.A(_08715_),
    .B(_08744_),
    .Y(_08745_));
 sky130_fd_sc_hd__xnor2_1 _16134_ (.A(_08713_),
    .B(_08745_),
    .Y(_08746_));
 sky130_fd_sc_hd__a21o_1 _16135_ (.A1(_08601_),
    .A2(_08610_),
    .B1(_08609_),
    .X(_08747_));
 sky130_fd_sc_hd__nand2_1 _16136_ (.A(_08616_),
    .B(_08622_),
    .Y(_08748_));
 sky130_fd_sc_hd__or4_1 _16137_ (.A(_07469_),
    .B(_08274_),
    .C(_08067_),
    .D(_07790_),
    .X(_08749_));
 sky130_fd_sc_hd__nand2_2 _16138_ (.A(_07384_),
    .B(_07385_),
    .Y(_08750_));
 sky130_fd_sc_hd__a2bb2o_1 _16139_ (.A1_N(_07469_),
    .A2_N(_08067_),
    .B1(_07520_),
    .B2(_08750_),
    .X(_08751_));
 sky130_fd_sc_hd__nand2_1 _16140_ (.A(_08749_),
    .B(_08751_),
    .Y(_08752_));
 sky130_fd_sc_hd__nor2_1 _16141_ (.A(_08596_),
    .B(_07886_),
    .Y(_08753_));
 sky130_fd_sc_hd__xnor2_1 _16142_ (.A(_08752_),
    .B(_08753_),
    .Y(_08754_));
 sky130_fd_sc_hd__or3_1 _16143_ (.A(_07800_),
    .B(_07712_),
    .C(_08603_),
    .X(_08755_));
 sky130_fd_sc_hd__o22ai_1 _16144_ (.A1(_08240_),
    .A2(_07712_),
    .B1(_07736_),
    .B2(_08241_),
    .Y(_08756_));
 sky130_fd_sc_hd__nand2_1 _16145_ (.A(_08755_),
    .B(_08756_),
    .Y(_08757_));
 sky130_fd_sc_hd__or2_1 _16146_ (.A(_07742_),
    .B(_07805_),
    .X(_08758_));
 sky130_fd_sc_hd__xnor2_1 _16147_ (.A(_08757_),
    .B(_08758_),
    .Y(_08759_));
 sky130_fd_sc_hd__clkbuf_4 _16148_ (.A(_07805_),
    .X(_08760_));
 sky130_fd_sc_hd__o31a_1 _16149_ (.A1(_07469_),
    .A2(_08760_),
    .A3(_08605_),
    .B1(_08602_),
    .X(_08761_));
 sky130_fd_sc_hd__xor2_1 _16150_ (.A(_08759_),
    .B(_08761_),
    .X(_08762_));
 sky130_fd_sc_hd__xnor2_1 _16151_ (.A(_08754_),
    .B(_08762_),
    .Y(_08763_));
 sky130_fd_sc_hd__a21o_1 _16152_ (.A1(_08748_),
    .A2(_08624_),
    .B1(_08763_),
    .X(_08764_));
 sky130_fd_sc_hd__nand3_1 _16153_ (.A(_08748_),
    .B(_08624_),
    .C(_08763_),
    .Y(_08765_));
 sky130_fd_sc_hd__nand2_1 _16154_ (.A(_08764_),
    .B(_08765_),
    .Y(_08766_));
 sky130_fd_sc_hd__xnor2_1 _16155_ (.A(_08747_),
    .B(_08766_),
    .Y(_08767_));
 sky130_fd_sc_hd__nand2_1 _16156_ (.A(_08619_),
    .B(_08618_),
    .Y(_08768_));
 sky130_fd_sc_hd__a22o_1 _16157_ (.A1(_08463_),
    .A2(_08617_),
    .B1(_08768_),
    .B2(_08621_),
    .X(_08769_));
 sky130_fd_sc_hd__a21boi_1 _16158_ (.A1(_08627_),
    .A2(_08637_),
    .B1_N(_08635_),
    .Y(_08770_));
 sky130_fd_sc_hd__clkbuf_4 _16159_ (.A(_07964_),
    .X(_08771_));
 sky130_fd_sc_hd__nand2_1 _16160_ (.A(_08771_),
    .B(_07837_),
    .Y(_08772_));
 sky130_fd_sc_hd__a21o_1 _16161_ (.A1(_08046_),
    .A2(_07837_),
    .B1(_08617_),
    .X(_08773_));
 sky130_fd_sc_hd__o21a_1 _16162_ (.A1(_08618_),
    .A2(_08772_),
    .B1(_08773_),
    .X(_08774_));
 sky130_fd_sc_hd__nor2_1 _16163_ (.A(_07858_),
    .B(_07685_),
    .Y(_08775_));
 sky130_fd_sc_hd__xor2_1 _16164_ (.A(_08774_),
    .B(_08775_),
    .X(_08776_));
 sky130_fd_sc_hd__xnor2_1 _16165_ (.A(_08770_),
    .B(_08776_),
    .Y(_08777_));
 sky130_fd_sc_hd__xor2_1 _16166_ (.A(_08769_),
    .B(_08777_),
    .X(_08778_));
 sky130_fd_sc_hd__clkinv_2 _16167_ (.A(_07814_),
    .Y(_08779_));
 sky130_fd_sc_hd__and2_2 _16168_ (.A(_07696_),
    .B(_08640_),
    .X(_08780_));
 sky130_fd_sc_hd__nand2_1 _16169_ (.A(_08629_),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .Y(_08781_));
 sky130_fd_sc_hd__or3_1 _16170_ (.A(_07229_),
    .B(_07234_),
    .C(_08474_),
    .X(_08782_));
 sky130_fd_sc_hd__o21ai_1 _16171_ (.A1(_07229_),
    .A2(_08474_),
    .B1(_07234_),
    .Y(_08783_));
 sky130_fd_sc_hd__a31o_1 _16172_ (.A1(_04933_),
    .A2(_08782_),
    .A3(_08783_),
    .B1(_07822_),
    .X(_08784_));
 sky130_fd_sc_hd__a21o_1 _16173_ (.A1(_08781_),
    .A2(_08784_),
    .B1(_07519_),
    .X(_08785_));
 sky130_fd_sc_hd__or4_1 _16174_ (.A(_07826_),
    .B(_07471_),
    .C(_08780_),
    .D(_08785_),
    .X(_08786_));
 sky130_fd_sc_hd__clkbuf_4 _16175_ (.A(_08785_),
    .X(_08787_));
 sky130_fd_sc_hd__nand2_2 _16176_ (.A(_07696_),
    .B(_08640_),
    .Y(_08788_));
 sky130_fd_sc_hd__a2bb2o_1 _16177_ (.A1_N(_07471_),
    .A2_N(_08787_),
    .B1(_08788_),
    .B2(_07697_),
    .X(_08789_));
 sky130_fd_sc_hd__nand4_1 _16178_ (.A(_08779_),
    .B(_08636_),
    .C(_08786_),
    .D(_08789_),
    .Y(_08790_));
 sky130_fd_sc_hd__a22o_1 _16179_ (.A1(_08779_),
    .A2(_08636_),
    .B1(_08786_),
    .B2(_08789_),
    .X(_08791_));
 sky130_fd_sc_hd__and2_1 _16180_ (.A(_08790_),
    .B(_08791_),
    .X(_08792_));
 sky130_fd_sc_hd__nand2_2 _16181_ (.A(_04938_),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .Y(_08793_));
 sky130_fd_sc_hd__a21o_1 _16182_ (.A1(_07824_),
    .A2(_08793_),
    .B1(_07835_),
    .X(_08794_));
 sky130_fd_sc_hd__nor2_1 _16183_ (.A(_08335_),
    .B(_08645_),
    .Y(_08795_));
 sky130_fd_sc_hd__xnor2_1 _16184_ (.A(_08794_),
    .B(_08795_),
    .Y(_08796_));
 sky130_fd_sc_hd__nor2_1 _16185_ (.A(_07847_),
    .B(_08634_),
    .Y(_08797_));
 sky130_fd_sc_hd__xnor2_1 _16186_ (.A(_08796_),
    .B(_08797_),
    .Y(_08798_));
 sky130_fd_sc_hd__nand2_1 _16187_ (.A(_08641_),
    .B(_08642_),
    .Y(_08799_));
 sky130_fd_sc_hd__o31a_1 _16188_ (.A1(_07843_),
    .A2(_08645_),
    .A3(_08643_),
    .B1(_08799_),
    .X(_08800_));
 sky130_fd_sc_hd__xor2_1 _16189_ (.A(_08798_),
    .B(_08800_),
    .X(_08801_));
 sky130_fd_sc_hd__xnor2_1 _16190_ (.A(_08792_),
    .B(_08801_),
    .Y(_08802_));
 sky130_fd_sc_hd__nor2_1 _16191_ (.A(_08647_),
    .B(_08648_),
    .Y(_08803_));
 sky130_fd_sc_hd__a21oi_1 _16192_ (.A1(_08639_),
    .A2(_08649_),
    .B1(_08803_),
    .Y(_08804_));
 sky130_fd_sc_hd__xor2_1 _16193_ (.A(_08802_),
    .B(_08804_),
    .X(_08805_));
 sky130_fd_sc_hd__xnor2_1 _16194_ (.A(_08778_),
    .B(_08805_),
    .Y(_08806_));
 sky130_fd_sc_hd__nor2_1 _16195_ (.A(_08650_),
    .B(_08651_),
    .Y(_08807_));
 sky130_fd_sc_hd__a21oi_1 _16196_ (.A1(_08626_),
    .A2(_08652_),
    .B1(_08807_),
    .Y(_08808_));
 sky130_fd_sc_hd__xor2_1 _16197_ (.A(_08806_),
    .B(_08808_),
    .X(_08809_));
 sky130_fd_sc_hd__xnor2_1 _16198_ (.A(_08767_),
    .B(_08809_),
    .Y(_08810_));
 sky130_fd_sc_hd__nor2_1 _16199_ (.A(_08653_),
    .B(_08654_),
    .Y(_08811_));
 sky130_fd_sc_hd__a21oi_1 _16200_ (.A1(_08614_),
    .A2(_08655_),
    .B1(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__xor2_1 _16201_ (.A(_08810_),
    .B(_08812_),
    .X(_08813_));
 sky130_fd_sc_hd__xnor2_1 _16202_ (.A(_08746_),
    .B(_08813_),
    .Y(_08814_));
 sky130_fd_sc_hd__nor2_1 _16203_ (.A(_08656_),
    .B(_08657_),
    .Y(_08815_));
 sky130_fd_sc_hd__a21oi_1 _16204_ (.A1(_08658_),
    .A2(_08685_),
    .B1(_08815_),
    .Y(_08816_));
 sky130_fd_sc_hd__or2_1 _16205_ (.A(_08814_),
    .B(_08816_),
    .X(_08817_));
 sky130_fd_sc_hd__nand2_1 _16206_ (.A(_08814_),
    .B(_08816_),
    .Y(_08818_));
 sky130_fd_sc_hd__nand2_1 _16207_ (.A(_08817_),
    .B(_08818_),
    .Y(_08819_));
 sky130_fd_sc_hd__or2b_1 _16208_ (.A(_08684_),
    .B_N(_08659_),
    .X(_08820_));
 sky130_fd_sc_hd__a21boi_1 _16209_ (.A1(_08661_),
    .A2(_08683_),
    .B1_N(_08820_),
    .Y(_08821_));
 sky130_fd_sc_hd__xnor2_1 _16210_ (.A(_08819_),
    .B(_08821_),
    .Y(_08822_));
 sky130_fd_sc_hd__o21a_1 _16211_ (.A1(_08691_),
    .A2(_08692_),
    .B1(_08689_),
    .X(_08823_));
 sky130_fd_sc_hd__xor2_1 _16212_ (.A(_08822_),
    .B(_08823_),
    .X(_08824_));
 sky130_fd_sc_hd__nand2_1 _16213_ (.A(_08711_),
    .B(_08824_),
    .Y(_08825_));
 sky130_fd_sc_hd__or2_1 _16214_ (.A(_08711_),
    .B(_08824_),
    .X(_08826_));
 sky130_fd_sc_hd__and2_2 _16215_ (.A(_08825_),
    .B(_08826_),
    .X(_08827_));
 sky130_fd_sc_hd__xnor2_4 _16216_ (.A(_08710_),
    .B(_08827_),
    .Y(_08828_));
 sky130_fd_sc_hd__clkinv_2 _16217_ (.A(\rbzero.debug_overlay.playerY[-4] ),
    .Y(_08829_));
 sky130_fd_sc_hd__mux2_1 _16218_ (.A0(_08829_),
    .A1(_07410_),
    .S(_07343_),
    .X(_08830_));
 sky130_fd_sc_hd__nor2_1 _16219_ (.A(_08828_),
    .B(_08830_),
    .Y(_08831_));
 sky130_fd_sc_hd__and2_1 _16220_ (.A(_08828_),
    .B(_08830_),
    .X(_08832_));
 sky130_fd_sc_hd__nor2_1 _16221_ (.A(_08831_),
    .B(_08832_),
    .Y(_08833_));
 sky130_fd_sc_hd__o21ba_1 _16222_ (.A1(_08704_),
    .A2(_08705_),
    .B1_N(_08702_),
    .X(_08834_));
 sky130_fd_sc_hd__xnor2_1 _16223_ (.A(_08833_),
    .B(_08834_),
    .Y(_08835_));
 sky130_fd_sc_hd__xnor2_1 _16224_ (.A(_08585_),
    .B(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__nand2_1 _16225_ (.A(_07338_),
    .B(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__o211a_1 _16226_ (.A1(\rbzero.wall_tracer.texu[2] ),
    .A2(_07338_),
    .B1(_07266_),
    .C1(_08837_),
    .X(_00483_));
 sky130_fd_sc_hd__o21bai_1 _16227_ (.A1(_08832_),
    .A2(_08834_),
    .B1_N(_08831_),
    .Y(_08838_));
 sky130_fd_sc_hd__a21bo_1 _16228_ (.A1(_08710_),
    .A2(_08827_),
    .B1_N(_08825_),
    .X(_08839_));
 sky130_fd_sc_hd__or2_2 _16229_ (.A(_08822_),
    .B(_08823_),
    .X(_08840_));
 sky130_fd_sc_hd__or2b_1 _16230_ (.A(_08664_),
    .B_N(_08727_),
    .X(_08841_));
 sky130_fd_sc_hd__or2b_1 _16231_ (.A(_08745_),
    .B_N(_08713_),
    .X(_08842_));
 sky130_fd_sc_hd__a21boi_1 _16232_ (.A1(_08715_),
    .A2(_08744_),
    .B1_N(_08842_),
    .Y(_08843_));
 sky130_fd_sc_hd__nor2_2 _16233_ (.A(_08841_),
    .B(_08843_),
    .Y(_08844_));
 sky130_fd_sc_hd__and2_1 _16234_ (.A(_08841_),
    .B(_08843_),
    .X(_08845_));
 sky130_fd_sc_hd__nor2_1 _16235_ (.A(_08844_),
    .B(_08845_),
    .Y(_08846_));
 sky130_fd_sc_hd__a21o_1 _16236_ (.A1(_08728_),
    .A2(_08743_),
    .B1(_08741_),
    .X(_08847_));
 sky130_fd_sc_hd__or2b_1 _16237_ (.A(_08766_),
    .B_N(_08747_),
    .X(_08848_));
 sky130_fd_sc_hd__or3b_1 _16238_ (.A(_08629_),
    .B(_04939_),
    .C_N(\rbzero.wall_tracer.visualWallDist[9] ),
    .X(_08849_));
 sky130_fd_sc_hd__buf_2 _16239_ (.A(_08849_),
    .X(_08850_));
 sky130_fd_sc_hd__buf_2 _16240_ (.A(_08850_),
    .X(_08851_));
 sky130_fd_sc_hd__clkbuf_4 _16241_ (.A(_08851_),
    .X(_08852_));
 sky130_fd_sc_hd__or2_1 _16242_ (.A(_07625_),
    .B(_08852_),
    .X(_08853_));
 sky130_fd_sc_hd__or4b_1 _16243_ (.A(_07792_),
    .B(_07788_),
    .C(_08717_),
    .D_N(\rbzero.wall_tracer.visualWallDist[7] ),
    .X(_08854_));
 sky130_fd_sc_hd__nor2_2 _16244_ (.A(_04938_),
    .B(_08663_),
    .Y(_08855_));
 sky130_fd_sc_hd__a2bb2o_1 _16245_ (.A1_N(_07878_),
    .A2_N(_08718_),
    .B1(_08855_),
    .B2(_07521_),
    .X(_08856_));
 sky130_fd_sc_hd__nand2_1 _16246_ (.A(_08854_),
    .B(_08856_),
    .Y(_08857_));
 sky130_fd_sc_hd__or2_1 _16247_ (.A(_08429_),
    .B(_08724_),
    .X(_08858_));
 sky130_fd_sc_hd__xnor2_1 _16248_ (.A(_08857_),
    .B(_08858_),
    .Y(_08859_));
 sky130_fd_sc_hd__o31a_1 _16249_ (.A1(_07625_),
    .A2(_08721_),
    .A3(_08725_),
    .B1(_08719_),
    .X(_08860_));
 sky130_fd_sc_hd__xor2_1 _16250_ (.A(_08859_),
    .B(_08860_),
    .X(_08861_));
 sky130_fd_sc_hd__xnor2_1 _16251_ (.A(_08853_),
    .B(_08861_),
    .Y(_08862_));
 sky130_fd_sc_hd__a21bo_1 _16252_ (.A1(_08733_),
    .A2(_08736_),
    .B1_N(_08731_),
    .X(_08863_));
 sky130_fd_sc_hd__a21bo_1 _16253_ (.A1(_08751_),
    .A2(_08753_),
    .B1_N(_08749_),
    .X(_08864_));
 sky130_fd_sc_hd__or4b_1 _16254_ (.A(_08592_),
    .B(_08296_),
    .C(_07621_),
    .D_N(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_08865_));
 sky130_fd_sc_hd__a2bb2o_1 _16255_ (.A1_N(_08592_),
    .A2_N(_08732_),
    .B1(_08536_),
    .B2(_08507_),
    .X(_08866_));
 sky130_fd_sc_hd__nand2_1 _16256_ (.A(_08865_),
    .B(_08866_),
    .Y(_08867_));
 sky130_fd_sc_hd__nor2_1 _16257_ (.A(_08510_),
    .B(_08735_),
    .Y(_08868_));
 sky130_fd_sc_hd__xor2_1 _16258_ (.A(_08867_),
    .B(_08868_),
    .X(_08869_));
 sky130_fd_sc_hd__xnor2_1 _16259_ (.A(_08864_),
    .B(_08869_),
    .Y(_08870_));
 sky130_fd_sc_hd__xnor2_1 _16260_ (.A(_08863_),
    .B(_08870_),
    .Y(_08871_));
 sky130_fd_sc_hd__and2b_1 _16261_ (.A_N(_08737_),
    .B(_08730_),
    .X(_08872_));
 sky130_fd_sc_hd__a21oi_1 _16262_ (.A1(_08729_),
    .A2(_08738_),
    .B1(_08872_),
    .Y(_08873_));
 sky130_fd_sc_hd__nor2_1 _16263_ (.A(_08871_),
    .B(_08873_),
    .Y(_08874_));
 sky130_fd_sc_hd__and2_1 _16264_ (.A(_08871_),
    .B(_08873_),
    .X(_08875_));
 sky130_fd_sc_hd__nor2_1 _16265_ (.A(_08874_),
    .B(_08875_),
    .Y(_08876_));
 sky130_fd_sc_hd__xnor2_1 _16266_ (.A(_08862_),
    .B(_08876_),
    .Y(_08877_));
 sky130_fd_sc_hd__a21o_1 _16267_ (.A1(_08764_),
    .A2(_08848_),
    .B1(_08877_),
    .X(_08878_));
 sky130_fd_sc_hd__nand3_1 _16268_ (.A(_08764_),
    .B(_08848_),
    .C(_08877_),
    .Y(_08879_));
 sky130_fd_sc_hd__nand2_1 _16269_ (.A(_08878_),
    .B(_08879_),
    .Y(_08880_));
 sky130_fd_sc_hd__xnor2_1 _16270_ (.A(_08847_),
    .B(_08880_),
    .Y(_08881_));
 sky130_fd_sc_hd__nor2_1 _16271_ (.A(_08759_),
    .B(_08761_),
    .Y(_08882_));
 sky130_fd_sc_hd__a21o_1 _16272_ (.A1(_08754_),
    .A2(_08762_),
    .B1(_08882_),
    .X(_08883_));
 sky130_fd_sc_hd__and2b_1 _16273_ (.A_N(_08770_),
    .B(_08776_),
    .X(_08884_));
 sky130_fd_sc_hd__a21o_1 _16274_ (.A1(_08769_),
    .A2(_08777_),
    .B1(_08884_),
    .X(_08885_));
 sky130_fd_sc_hd__or4_1 _16275_ (.A(_07742_),
    .B(_08223_),
    .C(_07591_),
    .D(_07790_),
    .X(_08886_));
 sky130_fd_sc_hd__a2bb2o_1 _16276_ (.A1_N(_07742_),
    .A2_N(_07591_),
    .B1(_07520_),
    .B2(_08135_),
    .X(_08887_));
 sky130_fd_sc_hd__nand2_1 _16277_ (.A(_08886_),
    .B(_08887_),
    .Y(_08888_));
 sky130_fd_sc_hd__or3_1 _16278_ (.A(_08274_),
    .B(_07598_),
    .C(_08888_),
    .X(_08889_));
 sky130_fd_sc_hd__buf_2 _16279_ (.A(_08274_),
    .X(_08890_));
 sky130_fd_sc_hd__o21ai_1 _16280_ (.A1(_08890_),
    .A2(_07886_),
    .B1(_08888_),
    .Y(_08891_));
 sky130_fd_sc_hd__and2_1 _16281_ (.A(_08889_),
    .B(_08891_),
    .X(_08892_));
 sky130_fd_sc_hd__nand2_1 _16282_ (.A(_07672_),
    .B(_07673_),
    .Y(_08893_));
 sky130_fd_sc_hd__and4b_1 _16283_ (.A_N(_07890_),
    .B(_07553_),
    .C(_08893_),
    .D(_07726_),
    .X(_08894_));
 sky130_fd_sc_hd__o22a_1 _16284_ (.A1(_08240_),
    .A2(_07685_),
    .B1(_07712_),
    .B2(_07800_),
    .X(_08895_));
 sky130_fd_sc_hd__nor2_1 _16285_ (.A(_08894_),
    .B(_08895_),
    .Y(_08896_));
 sky130_fd_sc_hd__nor2_1 _16286_ (.A(_08760_),
    .B(_07736_),
    .Y(_08897_));
 sky130_fd_sc_hd__xnor2_2 _16287_ (.A(_08896_),
    .B(_08897_),
    .Y(_08898_));
 sky130_fd_sc_hd__o31a_1 _16288_ (.A1(_07742_),
    .A2(_08760_),
    .A3(_08757_),
    .B1(_08755_),
    .X(_08899_));
 sky130_fd_sc_hd__xor2_2 _16289_ (.A(_08898_),
    .B(_08899_),
    .X(_08900_));
 sky130_fd_sc_hd__xor2_2 _16290_ (.A(_08892_),
    .B(_08900_),
    .X(_08901_));
 sky130_fd_sc_hd__xnor2_1 _16291_ (.A(_08885_),
    .B(_08901_),
    .Y(_08902_));
 sky130_fd_sc_hd__xnor2_1 _16292_ (.A(_08883_),
    .B(_08902_),
    .Y(_08903_));
 sky130_fd_sc_hd__a2bb2o_1 _16293_ (.A1_N(_08618_),
    .A2_N(_08772_),
    .B1(_08773_),
    .B2(_08775_),
    .X(_08904_));
 sky130_fd_sc_hd__nand2_1 _16294_ (.A(_08046_),
    .B(_08636_),
    .Y(_08905_));
 sky130_fd_sc_hd__and4_1 _16295_ (.A(_08046_),
    .B(_08771_),
    .C(_07837_),
    .D(_08636_),
    .X(_08906_));
 sky130_fd_sc_hd__a21oi_1 _16296_ (.A1(_08772_),
    .A2(_08905_),
    .B1(_08906_),
    .Y(_08907_));
 sky130_fd_sc_hd__nor2_1 _16297_ (.A(_07858_),
    .B(_07817_),
    .Y(_08908_));
 sky130_fd_sc_hd__xnor2_1 _16298_ (.A(_08907_),
    .B(_08908_),
    .Y(_08909_));
 sky130_fd_sc_hd__a21o_1 _16299_ (.A1(_08786_),
    .A2(_08790_),
    .B1(_08909_),
    .X(_08910_));
 sky130_fd_sc_hd__nand3_1 _16300_ (.A(_08786_),
    .B(_08790_),
    .C(_08909_),
    .Y(_08911_));
 sky130_fd_sc_hd__and3_1 _16301_ (.A(_08904_),
    .B(_08910_),
    .C(_08911_),
    .X(_08912_));
 sky130_fd_sc_hd__a21oi_1 _16302_ (.A1(_08910_),
    .A2(_08911_),
    .B1(_08904_),
    .Y(_08913_));
 sky130_fd_sc_hd__nor2_1 _16303_ (.A(_08912_),
    .B(_08913_),
    .Y(_08914_));
 sky130_fd_sc_hd__nand2_1 _16304_ (.A(_08779_),
    .B(_08788_),
    .Y(_08915_));
 sky130_fd_sc_hd__and2_1 _16305_ (.A(_07824_),
    .B(_08793_),
    .X(_08916_));
 sky130_fd_sc_hd__clkbuf_4 _16306_ (.A(_08916_),
    .X(_08917_));
 sky130_fd_sc_hd__nand2_1 _16307_ (.A(_08629_),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .Y(_08918_));
 sky130_fd_sc_hd__nor4_2 _16308_ (.A(_07229_),
    .B(_07234_),
    .C(_07237_),
    .D(_08474_),
    .Y(_08919_));
 sky130_fd_sc_hd__o31a_1 _16309_ (.A1(_07229_),
    .A2(_07234_),
    .A3(_08474_),
    .B1(_07237_),
    .X(_08920_));
 sky130_fd_sc_hd__o31ai_4 _16310_ (.A1(_07338_),
    .A2(_08919_),
    .A3(_08920_),
    .B1(_07694_),
    .Y(_08921_));
 sky130_fd_sc_hd__a21o_1 _16311_ (.A1(_08918_),
    .A2(_08921_),
    .B1(_04938_),
    .X(_08922_));
 sky130_fd_sc_hd__clkbuf_4 _16312_ (.A(_08922_),
    .X(_08923_));
 sky130_fd_sc_hd__and4bb_1 _16313_ (.A_N(_08917_),
    .B_N(_08923_),
    .C(_07697_),
    .D(_07698_),
    .X(_08924_));
 sky130_fd_sc_hd__o22a_1 _16314_ (.A1(_07826_),
    .A2(_08917_),
    .B1(_08923_),
    .B2(_07471_),
    .X(_08925_));
 sky130_fd_sc_hd__nor2_1 _16315_ (.A(_08924_),
    .B(_08925_),
    .Y(_08926_));
 sky130_fd_sc_hd__xnor2_1 _16316_ (.A(_08915_),
    .B(_08926_),
    .Y(_08927_));
 sky130_fd_sc_hd__nand2_2 _16317_ (.A(_04937_),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .Y(_08928_));
 sky130_fd_sc_hd__a21oi_1 _16318_ (.A1(_08478_),
    .A2(_08928_),
    .B1(_07835_),
    .Y(_08929_));
 sky130_fd_sc_hd__and3_1 _16319_ (.A(_04929_),
    .B(_07652_),
    .C(_08633_),
    .X(_08930_));
 sky130_fd_sc_hd__xnor2_1 _16320_ (.A(_08929_),
    .B(_08930_),
    .Y(_08931_));
 sky130_fd_sc_hd__nor2_1 _16321_ (.A(_07847_),
    .B(_08787_),
    .Y(_08932_));
 sky130_fd_sc_hd__xnor2_1 _16322_ (.A(_08931_),
    .B(_08932_),
    .Y(_08933_));
 sky130_fd_sc_hd__and2b_1 _16323_ (.A_N(_08794_),
    .B(_08795_),
    .X(_08934_));
 sky130_fd_sc_hd__a21oi_1 _16324_ (.A1(_08796_),
    .A2(_08797_),
    .B1(_08934_),
    .Y(_08935_));
 sky130_fd_sc_hd__xnor2_1 _16325_ (.A(_08933_),
    .B(_08935_),
    .Y(_08936_));
 sky130_fd_sc_hd__xor2_1 _16326_ (.A(_08927_),
    .B(_08936_),
    .X(_08937_));
 sky130_fd_sc_hd__nor2_1 _16327_ (.A(_08798_),
    .B(_08800_),
    .Y(_08938_));
 sky130_fd_sc_hd__a21o_1 _16328_ (.A1(_08792_),
    .A2(_08801_),
    .B1(_08938_),
    .X(_08939_));
 sky130_fd_sc_hd__xor2_1 _16329_ (.A(_08937_),
    .B(_08939_),
    .X(_08940_));
 sky130_fd_sc_hd__xor2_1 _16330_ (.A(_08914_),
    .B(_08940_),
    .X(_08941_));
 sky130_fd_sc_hd__nor2_1 _16331_ (.A(_08802_),
    .B(_08804_),
    .Y(_08942_));
 sky130_fd_sc_hd__a21o_1 _16332_ (.A1(_08778_),
    .A2(_08805_),
    .B1(_08942_),
    .X(_08943_));
 sky130_fd_sc_hd__xor2_1 _16333_ (.A(_08941_),
    .B(_08943_),
    .X(_08944_));
 sky130_fd_sc_hd__xor2_1 _16334_ (.A(_08903_),
    .B(_08944_),
    .X(_08945_));
 sky130_fd_sc_hd__nor2_1 _16335_ (.A(_08806_),
    .B(_08808_),
    .Y(_08946_));
 sky130_fd_sc_hd__a21o_1 _16336_ (.A1(_08767_),
    .A2(_08809_),
    .B1(_08946_),
    .X(_08947_));
 sky130_fd_sc_hd__xor2_1 _16337_ (.A(_08945_),
    .B(_08947_),
    .X(_08948_));
 sky130_fd_sc_hd__xnor2_1 _16338_ (.A(_08881_),
    .B(_08948_),
    .Y(_08949_));
 sky130_fd_sc_hd__nor2_1 _16339_ (.A(_08810_),
    .B(_08812_),
    .Y(_08950_));
 sky130_fd_sc_hd__a21oi_1 _16340_ (.A1(_08746_),
    .A2(_08813_),
    .B1(_08950_),
    .Y(_08951_));
 sky130_fd_sc_hd__xor2_1 _16341_ (.A(_08949_),
    .B(_08951_),
    .X(_08952_));
 sky130_fd_sc_hd__xnor2_1 _16342_ (.A(_08846_),
    .B(_08952_),
    .Y(_08953_));
 sky130_fd_sc_hd__o21a_1 _16343_ (.A1(_08819_),
    .A2(_08821_),
    .B1(_08817_),
    .X(_08954_));
 sky130_fd_sc_hd__or2_2 _16344_ (.A(_08953_),
    .B(_08954_),
    .X(_08955_));
 sky130_fd_sc_hd__nand2_1 _16345_ (.A(_08953_),
    .B(_08954_),
    .Y(_08956_));
 sky130_fd_sc_hd__and2_2 _16346_ (.A(_08955_),
    .B(_08956_),
    .X(_08957_));
 sky130_fd_sc_hd__xnor2_4 _16347_ (.A(_08840_),
    .B(_08957_),
    .Y(_08958_));
 sky130_fd_sc_hd__xor2_4 _16348_ (.A(_08839_),
    .B(_08958_),
    .X(_08959_));
 sky130_fd_sc_hd__clkinv_2 _16349_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .Y(_08960_));
 sky130_fd_sc_hd__mux2_1 _16350_ (.A0(_08960_),
    .A1(_07537_),
    .S(_07343_),
    .X(_08961_));
 sky130_fd_sc_hd__xnor2_1 _16351_ (.A(_08959_),
    .B(_08961_),
    .Y(_08962_));
 sky130_fd_sc_hd__xnor2_1 _16352_ (.A(_08838_),
    .B(_08962_),
    .Y(_08963_));
 sky130_fd_sc_hd__and2_1 _16353_ (.A(_08585_),
    .B(_08963_),
    .X(_08964_));
 sky130_fd_sc_hd__nor2_1 _16354_ (.A(_08585_),
    .B(_08963_),
    .Y(_08965_));
 sky130_fd_sc_hd__or3_1 _16355_ (.A(_04933_),
    .B(_08964_),
    .C(_08965_),
    .X(_08966_));
 sky130_fd_sc_hd__o211a_1 _16356_ (.A1(\rbzero.wall_tracer.texu[3] ),
    .A2(_07338_),
    .B1(_07266_),
    .C1(_08966_),
    .X(_00484_));
 sky130_fd_sc_hd__and2b_1 _16357_ (.A_N(_08961_),
    .B(_08959_),
    .X(_08967_));
 sky130_fd_sc_hd__a21o_1 _16358_ (.A1(_08838_),
    .A2(_08962_),
    .B1(_08967_),
    .X(_08968_));
 sky130_fd_sc_hd__or2b_1 _16359_ (.A(_08880_),
    .B_N(_08847_),
    .X(_08969_));
 sky130_fd_sc_hd__or2b_1 _16360_ (.A(_08853_),
    .B_N(_08861_),
    .X(_08970_));
 sky130_fd_sc_hd__o21a_1 _16361_ (.A1(_08859_),
    .A2(_08860_),
    .B1(_08970_),
    .X(_08971_));
 sky130_fd_sc_hd__a21oi_2 _16362_ (.A1(_08878_),
    .A2(_08969_),
    .B1(_08971_),
    .Y(_08972_));
 sky130_fd_sc_hd__and3_1 _16363_ (.A(_08878_),
    .B(_08969_),
    .C(_08971_),
    .X(_08973_));
 sky130_fd_sc_hd__nor2_1 _16364_ (.A(_08972_),
    .B(_08973_),
    .Y(_08974_));
 sky130_fd_sc_hd__a21o_1 _16365_ (.A1(_08862_),
    .A2(_08876_),
    .B1(_08874_),
    .X(_08975_));
 sky130_fd_sc_hd__nand2_1 _16366_ (.A(_08885_),
    .B(_08901_),
    .Y(_08976_));
 sky130_fd_sc_hd__or2b_1 _16367_ (.A(_08902_),
    .B_N(_08883_),
    .X(_08977_));
 sky130_fd_sc_hd__or3_4 _16368_ (.A(_05301_),
    .B(_08629_),
    .C(_04939_),
    .X(_08978_));
 sky130_fd_sc_hd__clkbuf_4 _16369_ (.A(_08978_),
    .X(_08979_));
 sky130_fd_sc_hd__or2_1 _16370_ (.A(_07625_),
    .B(_08979_),
    .X(_08980_));
 sky130_fd_sc_hd__nor2_1 _16371_ (.A(_08429_),
    .B(_08852_),
    .Y(_08981_));
 sky130_fd_sc_hd__xnor2_1 _16372_ (.A(_08980_),
    .B(_08981_),
    .Y(_08982_));
 sky130_fd_sc_hd__nor2_1 _16373_ (.A(_07515_),
    .B(_08723_),
    .Y(_08983_));
 sky130_fd_sc_hd__or2_1 _16374_ (.A(_07519_),
    .B(_08663_),
    .X(_08984_));
 sky130_fd_sc_hd__buf_2 _16375_ (.A(_08984_),
    .X(_08985_));
 sky130_fd_sc_hd__o22a_1 _16376_ (.A1(_07880_),
    .A2(_08717_),
    .B1(_08985_),
    .B2(_07878_),
    .X(_08986_));
 sky130_fd_sc_hd__or4_1 _16377_ (.A(_07792_),
    .B(_07880_),
    .C(_08717_),
    .D(_08984_),
    .X(_08987_));
 sky130_fd_sc_hd__and2b_1 _16378_ (.A_N(_08986_),
    .B(_08987_),
    .X(_08988_));
 sky130_fd_sc_hd__xnor2_1 _16379_ (.A(_08983_),
    .B(_08988_),
    .Y(_08989_));
 sky130_fd_sc_hd__o31a_1 _16380_ (.A1(_08429_),
    .A2(_08724_),
    .A3(_08857_),
    .B1(_08854_),
    .X(_08990_));
 sky130_fd_sc_hd__nor2_1 _16381_ (.A(_08989_),
    .B(_08990_),
    .Y(_08991_));
 sky130_fd_sc_hd__and2_1 _16382_ (.A(_08989_),
    .B(_08990_),
    .X(_08992_));
 sky130_fd_sc_hd__nor2_1 _16383_ (.A(_08991_),
    .B(_08992_),
    .Y(_08993_));
 sky130_fd_sc_hd__xor2_1 _16384_ (.A(_08982_),
    .B(_08993_),
    .X(_08994_));
 sky130_fd_sc_hd__a21bo_1 _16385_ (.A1(_08866_),
    .A2(_08868_),
    .B1_N(_08865_),
    .X(_08995_));
 sky130_fd_sc_hd__nand2_1 _16386_ (.A(_08886_),
    .B(_08889_),
    .Y(_08996_));
 sky130_fd_sc_hd__nor2_1 _16387_ (.A(_08599_),
    .B(_07916_),
    .Y(_08997_));
 sky130_fd_sc_hd__o22a_1 _16388_ (.A1(_08274_),
    .A2(_07621_),
    .B1(_08671_),
    .B2(_08592_),
    .X(_08998_));
 sky130_fd_sc_hd__or4_1 _16389_ (.A(_08274_),
    .B(_08592_),
    .C(_07620_),
    .D(_08671_),
    .X(_08999_));
 sky130_fd_sc_hd__and2b_1 _16390_ (.A_N(_08998_),
    .B(_08999_),
    .X(_09000_));
 sky130_fd_sc_hd__xnor2_1 _16391_ (.A(_08997_),
    .B(_09000_),
    .Y(_09001_));
 sky130_fd_sc_hd__xnor2_1 _16392_ (.A(_08996_),
    .B(_09001_),
    .Y(_09002_));
 sky130_fd_sc_hd__xnor2_1 _16393_ (.A(_08995_),
    .B(_09002_),
    .Y(_09003_));
 sky130_fd_sc_hd__and2b_1 _16394_ (.A_N(_08869_),
    .B(_08864_),
    .X(_09004_));
 sky130_fd_sc_hd__a21oi_1 _16395_ (.A1(_08863_),
    .A2(_08870_),
    .B1(_09004_),
    .Y(_09005_));
 sky130_fd_sc_hd__nor2_1 _16396_ (.A(_09003_),
    .B(_09005_),
    .Y(_09006_));
 sky130_fd_sc_hd__and2_1 _16397_ (.A(_09003_),
    .B(_09005_),
    .X(_09007_));
 sky130_fd_sc_hd__nor2_1 _16398_ (.A(_09006_),
    .B(_09007_),
    .Y(_09008_));
 sky130_fd_sc_hd__xnor2_1 _16399_ (.A(_08994_),
    .B(_09008_),
    .Y(_09009_));
 sky130_fd_sc_hd__a21o_1 _16400_ (.A1(_08976_),
    .A2(_08977_),
    .B1(_09009_),
    .X(_09010_));
 sky130_fd_sc_hd__nand3_1 _16401_ (.A(_08976_),
    .B(_08977_),
    .C(_09009_),
    .Y(_09011_));
 sky130_fd_sc_hd__nand2_1 _16402_ (.A(_09010_),
    .B(_09011_),
    .Y(_09012_));
 sky130_fd_sc_hd__xnor2_1 _16403_ (.A(_08975_),
    .B(_09012_),
    .Y(_09013_));
 sky130_fd_sc_hd__nor2_1 _16404_ (.A(_08898_),
    .B(_08899_),
    .Y(_09014_));
 sky130_fd_sc_hd__a21o_1 _16405_ (.A1(_08892_),
    .A2(_08900_),
    .B1(_09014_),
    .X(_09015_));
 sky130_fd_sc_hd__a21bo_1 _16406_ (.A1(_08904_),
    .A2(_08911_),
    .B1_N(_08910_),
    .X(_09016_));
 sky130_fd_sc_hd__or4_1 _16407_ (.A(_08086_),
    .B(_07591_),
    .C(_07790_),
    .D(_07735_),
    .X(_09017_));
 sky130_fd_sc_hd__nand2_2 _16408_ (.A(_07439_),
    .B(_07440_),
    .Y(_09018_));
 sky130_fd_sc_hd__a2bb2o_1 _16409_ (.A1_N(_07591_),
    .A2_N(_07736_),
    .B1(_07520_),
    .B2(_09018_),
    .X(_09019_));
 sky130_fd_sc_hd__nand2_1 _16410_ (.A(_09017_),
    .B(_09019_),
    .Y(_09020_));
 sky130_fd_sc_hd__or3_1 _16411_ (.A(_08223_),
    .B(_07598_),
    .C(_09020_),
    .X(_09021_));
 sky130_fd_sc_hd__buf_2 _16412_ (.A(_08223_),
    .X(_09022_));
 sky130_fd_sc_hd__o21ai_1 _16413_ (.A1(_09022_),
    .A2(_07886_),
    .B1(_09020_),
    .Y(_09023_));
 sky130_fd_sc_hd__and2_1 _16414_ (.A(_09021_),
    .B(_09023_),
    .X(_09024_));
 sky130_fd_sc_hd__or4_1 _16415_ (.A(_07890_),
    .B(_07800_),
    .C(_07685_),
    .D(_07817_),
    .X(_09025_));
 sky130_fd_sc_hd__a2bb2o_1 _16416_ (.A1_N(_07890_),
    .A2_N(_07817_),
    .B1(_07553_),
    .B2(_08893_),
    .X(_09026_));
 sky130_fd_sc_hd__nand2_1 _16417_ (.A(_09025_),
    .B(_09026_),
    .Y(_09027_));
 sky130_fd_sc_hd__nor2_1 _16418_ (.A(_07567_),
    .B(_07712_),
    .Y(_09028_));
 sky130_fd_sc_hd__xor2_1 _16419_ (.A(_09027_),
    .B(_09028_),
    .X(_09029_));
 sky130_fd_sc_hd__a21oi_1 _16420_ (.A1(_08896_),
    .A2(_08897_),
    .B1(_08894_),
    .Y(_09030_));
 sky130_fd_sc_hd__xor2_1 _16421_ (.A(_09029_),
    .B(_09030_),
    .X(_09031_));
 sky130_fd_sc_hd__xnor2_1 _16422_ (.A(_09024_),
    .B(_09031_),
    .Y(_09032_));
 sky130_fd_sc_hd__xor2_1 _16423_ (.A(_09016_),
    .B(_09032_),
    .X(_09033_));
 sky130_fd_sc_hd__xnor2_1 _16424_ (.A(_09015_),
    .B(_09033_),
    .Y(_09034_));
 sky130_fd_sc_hd__a21o_1 _16425_ (.A1(_08907_),
    .A2(_08908_),
    .B1(_08906_),
    .X(_09035_));
 sky130_fd_sc_hd__o21bai_1 _16426_ (.A1(_08915_),
    .A2(_08925_),
    .B1_N(_08924_),
    .Y(_09036_));
 sky130_fd_sc_hd__and2_1 _16427_ (.A(_08046_),
    .B(_08636_),
    .X(_09037_));
 sky130_fd_sc_hd__a21o_1 _16428_ (.A1(_07696_),
    .A2(_08640_),
    .B1(_08272_),
    .X(_09038_));
 sky130_fd_sc_hd__nand2_1 _16429_ (.A(_08771_),
    .B(_08636_),
    .Y(_09039_));
 sky130_fd_sc_hd__a32o_1 _16430_ (.A1(_08771_),
    .A2(_08788_),
    .A3(_09037_),
    .B1(_09038_),
    .B2(_09039_),
    .X(_09040_));
 sky130_fd_sc_hd__nor2_1 _16431_ (.A(_07751_),
    .B(_07834_),
    .Y(_09041_));
 sky130_fd_sc_hd__xnor2_1 _16432_ (.A(_09040_),
    .B(_09041_),
    .Y(_09042_));
 sky130_fd_sc_hd__nand2_1 _16433_ (.A(_09036_),
    .B(_09042_),
    .Y(_09043_));
 sky130_fd_sc_hd__or2_1 _16434_ (.A(_09036_),
    .B(_09042_),
    .X(_09044_));
 sky130_fd_sc_hd__nand2_1 _16435_ (.A(_09043_),
    .B(_09044_),
    .Y(_09045_));
 sky130_fd_sc_hd__xnor2_1 _16436_ (.A(_09035_),
    .B(_09045_),
    .Y(_09046_));
 sky130_fd_sc_hd__a21o_1 _16437_ (.A1(_07824_),
    .A2(_08793_),
    .B1(_07468_),
    .X(_09047_));
 sky130_fd_sc_hd__a21o_1 _16438_ (.A1(_08478_),
    .A2(_08928_),
    .B1(_07826_),
    .X(_09048_));
 sky130_fd_sc_hd__o41a_1 _16439_ (.A1(_07229_),
    .A2(_07234_),
    .A3(_07237_),
    .A4(_08474_),
    .B1(_07241_),
    .X(_09049_));
 sky130_fd_sc_hd__a211o_1 _16440_ (.A1(_07240_),
    .A2(_08919_),
    .B1(_09049_),
    .C1(_07338_),
    .X(_09050_));
 sky130_fd_sc_hd__a22oi_4 _16441_ (.A1(_08629_),
    .A2(\rbzero.wall_tracer.stepDistY[10] ),
    .B1(_07694_),
    .B2(_09050_),
    .Y(_09051_));
 sky130_fd_sc_hd__nor2_1 _16442_ (.A(_08398_),
    .B(_09051_),
    .Y(_09052_));
 sky130_fd_sc_hd__xnor2_1 _16443_ (.A(_09048_),
    .B(_09052_),
    .Y(_09053_));
 sky130_fd_sc_hd__xnor2_1 _16444_ (.A(_09047_),
    .B(_09053_),
    .Y(_09054_));
 sky130_fd_sc_hd__mux2_4 _16445_ (.A0(\rbzero.wall_tracer.stepDistX[7] ),
    .A1(_08633_),
    .S(_04929_),
    .X(_09055_));
 sky130_fd_sc_hd__or4b_1 _16446_ (.A(_07835_),
    .B(_07680_),
    .C(_08785_),
    .D_N(_09055_),
    .X(_09056_));
 sky130_fd_sc_hd__a2bb2o_1 _16447_ (.A1_N(_07680_),
    .A2_N(_08787_),
    .B1(_09055_),
    .B2(_07838_),
    .X(_09057_));
 sky130_fd_sc_hd__nor2_1 _16448_ (.A(_07847_),
    .B(_08923_),
    .Y(_09058_));
 sky130_fd_sc_hd__nand3_1 _16449_ (.A(_09056_),
    .B(_09057_),
    .C(_09058_),
    .Y(_09059_));
 sky130_fd_sc_hd__a21o_1 _16450_ (.A1(_09056_),
    .A2(_09057_),
    .B1(_09058_),
    .X(_09060_));
 sky130_fd_sc_hd__nand2_1 _16451_ (.A(_08929_),
    .B(_08930_),
    .Y(_09061_));
 sky130_fd_sc_hd__o31ai_1 _16452_ (.A1(_07847_),
    .A2(_08787_),
    .A3(_08931_),
    .B1(_09061_),
    .Y(_09062_));
 sky130_fd_sc_hd__nand3_1 _16453_ (.A(_09059_),
    .B(_09060_),
    .C(_09062_),
    .Y(_09063_));
 sky130_fd_sc_hd__a21o_1 _16454_ (.A1(_09059_),
    .A2(_09060_),
    .B1(_09062_),
    .X(_09064_));
 sky130_fd_sc_hd__nand3_1 _16455_ (.A(_09054_),
    .B(_09063_),
    .C(_09064_),
    .Y(_09065_));
 sky130_fd_sc_hd__a21o_1 _16456_ (.A1(_09063_),
    .A2(_09064_),
    .B1(_09054_),
    .X(_09066_));
 sky130_fd_sc_hd__and2b_1 _16457_ (.A_N(_08935_),
    .B(_08933_),
    .X(_09067_));
 sky130_fd_sc_hd__a21o_1 _16458_ (.A1(_08927_),
    .A2(_08936_),
    .B1(_09067_),
    .X(_09068_));
 sky130_fd_sc_hd__nand3_1 _16459_ (.A(_09065_),
    .B(_09066_),
    .C(_09068_),
    .Y(_09069_));
 sky130_fd_sc_hd__a21o_1 _16460_ (.A1(_09065_),
    .A2(_09066_),
    .B1(_09068_),
    .X(_09070_));
 sky130_fd_sc_hd__nand3_1 _16461_ (.A(_09046_),
    .B(_09069_),
    .C(_09070_),
    .Y(_09071_));
 sky130_fd_sc_hd__a21o_1 _16462_ (.A1(_09069_),
    .A2(_09070_),
    .B1(_09046_),
    .X(_09072_));
 sky130_fd_sc_hd__nand2_1 _16463_ (.A(_08937_),
    .B(_08939_),
    .Y(_09073_));
 sky130_fd_sc_hd__a21bo_1 _16464_ (.A1(_08914_),
    .A2(_08940_),
    .B1_N(_09073_),
    .X(_09074_));
 sky130_fd_sc_hd__nand3_1 _16465_ (.A(_09071_),
    .B(_09072_),
    .C(_09074_),
    .Y(_09075_));
 sky130_fd_sc_hd__a21o_1 _16466_ (.A1(_09071_),
    .A2(_09072_),
    .B1(_09074_),
    .X(_09076_));
 sky130_fd_sc_hd__nand3_1 _16467_ (.A(_09034_),
    .B(_09075_),
    .C(_09076_),
    .Y(_09077_));
 sky130_fd_sc_hd__a21o_1 _16468_ (.A1(_09075_),
    .A2(_09076_),
    .B1(_09034_),
    .X(_09078_));
 sky130_fd_sc_hd__nand2_1 _16469_ (.A(_08941_),
    .B(_08943_),
    .Y(_09079_));
 sky130_fd_sc_hd__a21bo_1 _16470_ (.A1(_08903_),
    .A2(_08944_),
    .B1_N(_09079_),
    .X(_09080_));
 sky130_fd_sc_hd__nand3_1 _16471_ (.A(_09077_),
    .B(_09078_),
    .C(_09080_),
    .Y(_09081_));
 sky130_fd_sc_hd__a21o_1 _16472_ (.A1(_09077_),
    .A2(_09078_),
    .B1(_09080_),
    .X(_09082_));
 sky130_fd_sc_hd__nand3_1 _16473_ (.A(_09013_),
    .B(_09081_),
    .C(_09082_),
    .Y(_09083_));
 sky130_fd_sc_hd__a21o_1 _16474_ (.A1(_09081_),
    .A2(_09082_),
    .B1(_09013_),
    .X(_09084_));
 sky130_fd_sc_hd__nand2_1 _16475_ (.A(_08945_),
    .B(_08947_),
    .Y(_09085_));
 sky130_fd_sc_hd__a21bo_1 _16476_ (.A1(_08881_),
    .A2(_08948_),
    .B1_N(_09085_),
    .X(_09086_));
 sky130_fd_sc_hd__nand3_1 _16477_ (.A(_09083_),
    .B(_09084_),
    .C(_09086_),
    .Y(_09087_));
 sky130_fd_sc_hd__a21o_1 _16478_ (.A1(_09083_),
    .A2(_09084_),
    .B1(_09086_),
    .X(_09088_));
 sky130_fd_sc_hd__and3_1 _16479_ (.A(_08974_),
    .B(_09087_),
    .C(_09088_),
    .X(_09089_));
 sky130_fd_sc_hd__a21oi_1 _16480_ (.A1(_09087_),
    .A2(_09088_),
    .B1(_08974_),
    .Y(_09090_));
 sky130_fd_sc_hd__nor2_1 _16481_ (.A(_09089_),
    .B(_09090_),
    .Y(_09091_));
 sky130_fd_sc_hd__nor2_1 _16482_ (.A(_08949_),
    .B(_08951_),
    .Y(_09092_));
 sky130_fd_sc_hd__a21oi_1 _16483_ (.A1(_08846_),
    .A2(_08952_),
    .B1(_09092_),
    .Y(_09093_));
 sky130_fd_sc_hd__xnor2_1 _16484_ (.A(_09091_),
    .B(_09093_),
    .Y(_09094_));
 sky130_fd_sc_hd__xor2_2 _16485_ (.A(_08844_),
    .B(_09094_),
    .X(_09095_));
 sky130_fd_sc_hd__xor2_4 _16486_ (.A(_08955_),
    .B(_09095_),
    .X(_09096_));
 sky130_fd_sc_hd__nand2_1 _16487_ (.A(_08840_),
    .B(_08825_),
    .Y(_09097_));
 sky130_fd_sc_hd__a32oi_4 _16488_ (.A1(_08710_),
    .A2(_08827_),
    .A3(_08958_),
    .B1(_09097_),
    .B2(_08957_),
    .Y(_09098_));
 sky130_fd_sc_hd__xor2_4 _16489_ (.A(_09096_),
    .B(_09098_),
    .X(_09099_));
 sky130_fd_sc_hd__mux2_1 _16490_ (.A0(\rbzero.debug_overlay.playerY[-2] ),
    .A1(\rbzero.debug_overlay.playerX[-2] ),
    .S(_07343_),
    .X(_09100_));
 sky130_fd_sc_hd__or2_1 _16491_ (.A(_09099_),
    .B(_09100_),
    .X(_09101_));
 sky130_fd_sc_hd__nand2_1 _16492_ (.A(_09099_),
    .B(_09100_),
    .Y(_09102_));
 sky130_fd_sc_hd__nand2_1 _16493_ (.A(_09101_),
    .B(_09102_),
    .Y(_09103_));
 sky130_fd_sc_hd__xnor2_1 _16494_ (.A(_08585_),
    .B(_09103_),
    .Y(_09104_));
 sky130_fd_sc_hd__or2_1 _16495_ (.A(_08968_),
    .B(_09104_),
    .X(_09105_));
 sky130_fd_sc_hd__nand2_1 _16496_ (.A(_08968_),
    .B(_09104_),
    .Y(_09106_));
 sky130_fd_sc_hd__a21o_1 _16497_ (.A1(_09105_),
    .A2(_09106_),
    .B1(_04933_),
    .X(_09107_));
 sky130_fd_sc_hd__o211a_1 _16498_ (.A1(\rbzero.wall_tracer.texu[4] ),
    .A2(_07338_),
    .B1(_03819_),
    .C1(_09107_),
    .X(_00485_));
 sky130_fd_sc_hd__a21boi_1 _16499_ (.A1(_08968_),
    .A2(_09101_),
    .B1_N(_09102_),
    .Y(_09108_));
 sky130_fd_sc_hd__or2b_1 _16500_ (.A(_09012_),
    .B_N(_08975_),
    .X(_09109_));
 sky130_fd_sc_hd__or3_1 _16501_ (.A(_08429_),
    .B(_08852_),
    .C(_08980_),
    .X(_09110_));
 sky130_fd_sc_hd__xnor2_1 _16502_ (.A(_09110_),
    .B(_08991_),
    .Y(_09111_));
 sky130_fd_sc_hd__a21oi_1 _16503_ (.A1(_08982_),
    .A2(_08993_),
    .B1(_09111_),
    .Y(_09112_));
 sky130_fd_sc_hd__or3b_1 _16504_ (.A(_08629_),
    .B(_04938_),
    .C_N(\rbzero.wall_tracer.visualWallDist[11] ),
    .X(_09113_));
 sky130_fd_sc_hd__buf_2 _16505_ (.A(_09113_),
    .X(_09114_));
 sky130_fd_sc_hd__clkbuf_4 _16506_ (.A(_09114_),
    .X(_09115_));
 sky130_fd_sc_hd__or2_1 _16507_ (.A(_07632_),
    .B(_09115_),
    .X(_09116_));
 sky130_fd_sc_hd__xnor2_1 _16508_ (.A(_09112_),
    .B(_09116_),
    .Y(_09117_));
 sky130_fd_sc_hd__a21oi_1 _16509_ (.A1(_09010_),
    .A2(_09109_),
    .B1(_09117_),
    .Y(_09118_));
 sky130_fd_sc_hd__and3_1 _16510_ (.A(_09010_),
    .B(_09109_),
    .C(_09117_),
    .X(_09119_));
 sky130_fd_sc_hd__nor2_1 _16511_ (.A(_09118_),
    .B(_09119_),
    .Y(_09120_));
 sky130_fd_sc_hd__a21o_1 _16512_ (.A1(_08994_),
    .A2(_09008_),
    .B1(_09006_),
    .X(_09121_));
 sky130_fd_sc_hd__or2b_1 _16513_ (.A(_09032_),
    .B_N(_09016_),
    .X(_09122_));
 sky130_fd_sc_hd__or2b_1 _16514_ (.A(_09033_),
    .B_N(_09015_),
    .X(_09123_));
 sky130_fd_sc_hd__nor2_1 _16515_ (.A(_07878_),
    .B(_08723_),
    .Y(_09124_));
 sky130_fd_sc_hd__nor2_1 _16516_ (.A(_07515_),
    .B(_08850_),
    .Y(_09125_));
 sky130_fd_sc_hd__xnor2_1 _16517_ (.A(_09124_),
    .B(_09125_),
    .Y(_09126_));
 sky130_fd_sc_hd__nor2_1 _16518_ (.A(_08429_),
    .B(_08979_),
    .Y(_09127_));
 sky130_fd_sc_hd__xnor2_1 _16519_ (.A(_09126_),
    .B(_09127_),
    .Y(_09128_));
 sky130_fd_sc_hd__nor2_1 _16520_ (.A(_08510_),
    .B(_08985_),
    .Y(_09129_));
 sky130_fd_sc_hd__o22a_1 _16521_ (.A1(_08592_),
    .A2(_07916_),
    .B1(_08717_),
    .B2(_08296_),
    .X(_09130_));
 sky130_fd_sc_hd__or4_1 _16522_ (.A(_08592_),
    .B(_08296_),
    .C(_07916_),
    .D(_08716_),
    .X(_09131_));
 sky130_fd_sc_hd__and2b_1 _16523_ (.A_N(_09130_),
    .B(_09131_),
    .X(_09132_));
 sky130_fd_sc_hd__xnor2_1 _16524_ (.A(_09129_),
    .B(_09132_),
    .Y(_09133_));
 sky130_fd_sc_hd__o31a_1 _16525_ (.A1(_07515_),
    .A2(_08723_),
    .A3(_08986_),
    .B1(_08987_),
    .X(_09134_));
 sky130_fd_sc_hd__or2_1 _16526_ (.A(_09133_),
    .B(_09134_),
    .X(_09135_));
 sky130_fd_sc_hd__nand2_1 _16527_ (.A(_09133_),
    .B(_09134_),
    .Y(_09136_));
 sky130_fd_sc_hd__and2_1 _16528_ (.A(_09135_),
    .B(_09136_),
    .X(_09137_));
 sky130_fd_sc_hd__nand2_1 _16529_ (.A(_09128_),
    .B(_09137_),
    .Y(_09138_));
 sky130_fd_sc_hd__or2_1 _16530_ (.A(_09128_),
    .B(_09137_),
    .X(_09139_));
 sky130_fd_sc_hd__and2_1 _16531_ (.A(_09138_),
    .B(_09139_),
    .X(_09140_));
 sky130_fd_sc_hd__a21bo_1 _16532_ (.A1(_08997_),
    .A2(_09000_),
    .B1_N(_08999_),
    .X(_09141_));
 sky130_fd_sc_hd__nand2_1 _16533_ (.A(_09017_),
    .B(_09021_),
    .Y(_09142_));
 sky130_fd_sc_hd__nor2_1 _16534_ (.A(_08890_),
    .B(_08671_),
    .Y(_09143_));
 sky130_fd_sc_hd__o22a_1 _16535_ (.A1(_08086_),
    .A2(_07597_),
    .B1(_07621_),
    .B2(_08223_),
    .X(_09144_));
 sky130_fd_sc_hd__or4_1 _16536_ (.A(_08086_),
    .B(_08223_),
    .C(_07597_),
    .D(_07620_),
    .X(_09145_));
 sky130_fd_sc_hd__and2b_1 _16537_ (.A_N(_09144_),
    .B(_09145_),
    .X(_09146_));
 sky130_fd_sc_hd__xnor2_1 _16538_ (.A(_09143_),
    .B(_09146_),
    .Y(_09147_));
 sky130_fd_sc_hd__xnor2_1 _16539_ (.A(_09142_),
    .B(_09147_),
    .Y(_09148_));
 sky130_fd_sc_hd__xnor2_1 _16540_ (.A(_09141_),
    .B(_09148_),
    .Y(_09149_));
 sky130_fd_sc_hd__a21oi_1 _16541_ (.A1(_08886_),
    .A2(_08889_),
    .B1(_09001_),
    .Y(_09150_));
 sky130_fd_sc_hd__a21oi_1 _16542_ (.A1(_08995_),
    .A2(_09002_),
    .B1(_09150_),
    .Y(_09151_));
 sky130_fd_sc_hd__nor2_1 _16543_ (.A(_09149_),
    .B(_09151_),
    .Y(_09152_));
 sky130_fd_sc_hd__and2_1 _16544_ (.A(_09149_),
    .B(_09151_),
    .X(_09153_));
 sky130_fd_sc_hd__nor2_1 _16545_ (.A(_09152_),
    .B(_09153_),
    .Y(_09154_));
 sky130_fd_sc_hd__xnor2_1 _16546_ (.A(_09140_),
    .B(_09154_),
    .Y(_09155_));
 sky130_fd_sc_hd__a21o_1 _16547_ (.A1(_09122_),
    .A2(_09123_),
    .B1(_09155_),
    .X(_09156_));
 sky130_fd_sc_hd__nand3_1 _16548_ (.A(_09122_),
    .B(_09123_),
    .C(_09155_),
    .Y(_09157_));
 sky130_fd_sc_hd__nand2_1 _16549_ (.A(_09156_),
    .B(_09157_),
    .Y(_09158_));
 sky130_fd_sc_hd__xnor2_1 _16550_ (.A(_09121_),
    .B(_09158_),
    .Y(_09159_));
 sky130_fd_sc_hd__nor2_1 _16551_ (.A(_09029_),
    .B(_09030_),
    .Y(_09160_));
 sky130_fd_sc_hd__a21o_1 _16552_ (.A1(_09024_),
    .A2(_09031_),
    .B1(_09160_),
    .X(_09161_));
 sky130_fd_sc_hd__a21bo_1 _16553_ (.A1(_09035_),
    .A2(_09044_),
    .B1_N(_09043_),
    .X(_09162_));
 sky130_fd_sc_hd__buf_2 _16554_ (.A(_07793_),
    .X(_09163_));
 sky130_fd_sc_hd__o22a_1 _16555_ (.A1(_07805_),
    .A2(_07685_),
    .B1(_07712_),
    .B2(_08067_),
    .X(_09164_));
 sky130_fd_sc_hd__a31o_1 _16556_ (.A1(_09163_),
    .A2(_08893_),
    .A3(_09028_),
    .B1(_09164_),
    .X(_09165_));
 sky130_fd_sc_hd__buf_2 _16557_ (.A(_07936_),
    .X(_09166_));
 sky130_fd_sc_hd__nor2_1 _16558_ (.A(_08595_),
    .B(_09166_),
    .Y(_09167_));
 sky130_fd_sc_hd__xnor2_1 _16559_ (.A(_09165_),
    .B(_09167_),
    .Y(_09168_));
 sky130_fd_sc_hd__nor2_1 _16560_ (.A(_08241_),
    .B(_07817_),
    .Y(_09169_));
 sky130_fd_sc_hd__or2b_1 _16561_ (.A(_07890_),
    .B_N(_08636_),
    .X(_09170_));
 sky130_fd_sc_hd__and2b_1 _16562_ (.A_N(_07751_),
    .B(_08636_),
    .X(_09171_));
 sky130_fd_sc_hd__nor2_1 _16563_ (.A(_07890_),
    .B(_07834_),
    .Y(_09172_));
 sky130_fd_sc_hd__o32a_1 _16564_ (.A1(_07751_),
    .A2(_07834_),
    .A3(_09170_),
    .B1(_09171_),
    .B2(_09172_),
    .X(_09173_));
 sky130_fd_sc_hd__xnor2_1 _16565_ (.A(_09169_),
    .B(_09173_),
    .Y(_09174_));
 sky130_fd_sc_hd__o31a_1 _16566_ (.A1(_08760_),
    .A2(_07712_),
    .A3(_09027_),
    .B1(_09025_),
    .X(_09175_));
 sky130_fd_sc_hd__xor2_1 _16567_ (.A(_09174_),
    .B(_09175_),
    .X(_09176_));
 sky130_fd_sc_hd__xnor2_1 _16568_ (.A(_09168_),
    .B(_09176_),
    .Y(_09177_));
 sky130_fd_sc_hd__xnor2_1 _16569_ (.A(_09162_),
    .B(_09177_),
    .Y(_09178_));
 sky130_fd_sc_hd__and2_1 _16570_ (.A(_09161_),
    .B(_09178_),
    .X(_09179_));
 sky130_fd_sc_hd__nor2_1 _16571_ (.A(_09161_),
    .B(_09178_),
    .Y(_09180_));
 sky130_fd_sc_hd__nor2_1 _16572_ (.A(_09179_),
    .B(_09180_),
    .Y(_09181_));
 sky130_fd_sc_hd__clkbuf_4 _16573_ (.A(_07858_),
    .X(_09182_));
 sky130_fd_sc_hd__nand2_1 _16574_ (.A(_08771_),
    .B(_08788_),
    .Y(_09183_));
 sky130_fd_sc_hd__o32ai_2 _16575_ (.A1(_09182_),
    .A2(_07834_),
    .A3(_09040_),
    .B1(_09183_),
    .B2(_08905_),
    .Y(_09184_));
 sky130_fd_sc_hd__o21a_1 _16576_ (.A1(_08398_),
    .A2(_09051_),
    .B1(_09048_),
    .X(_09185_));
 sky130_fd_sc_hd__or3_1 _16577_ (.A(_08398_),
    .B(_09048_),
    .C(_09051_),
    .X(_09186_));
 sky130_fd_sc_hd__o21a_1 _16578_ (.A1(_09047_),
    .A2(_09185_),
    .B1(_09186_),
    .X(_09187_));
 sky130_fd_sc_hd__a21o_1 _16579_ (.A1(_08478_),
    .A2(_08928_),
    .B1(_08272_),
    .X(_09188_));
 sky130_fd_sc_hd__a21oi_1 _16580_ (.A1(_08478_),
    .A2(_08928_),
    .B1(_07814_),
    .Y(_09189_));
 sky130_fd_sc_hd__a21oi_1 _16581_ (.A1(_07824_),
    .A2(_08793_),
    .B1(_08272_),
    .Y(_09190_));
 sky130_fd_sc_hd__o22a_1 _16582_ (.A1(_09047_),
    .A2(_09188_),
    .B1(_09189_),
    .B2(_09190_),
    .X(_09191_));
 sky130_fd_sc_hd__xnor2_1 _16583_ (.A(_09183_),
    .B(_09191_),
    .Y(_09192_));
 sky130_fd_sc_hd__xnor2_1 _16584_ (.A(_09187_),
    .B(_09192_),
    .Y(_09193_));
 sky130_fd_sc_hd__nand2_1 _16585_ (.A(_09184_),
    .B(_09193_),
    .Y(_09194_));
 sky130_fd_sc_hd__or2_1 _16586_ (.A(_09184_),
    .B(_09193_),
    .X(_09195_));
 sky130_fd_sc_hd__and2_1 _16587_ (.A(_09194_),
    .B(_09195_),
    .X(_09196_));
 sky130_fd_sc_hd__a21boi_4 _16588_ (.A1(_04939_),
    .A2(\rbzero.wall_tracer.stepDistX[7] ),
    .B1_N(_08634_),
    .Y(_09197_));
 sky130_fd_sc_hd__inv_2 _16589_ (.A(_07243_),
    .Y(_09198_));
 sky130_fd_sc_hd__a31o_1 _16590_ (.A1(_07240_),
    .A2(_09198_),
    .A3(_08919_),
    .B1(_07337_),
    .X(_09199_));
 sky130_fd_sc_hd__a22oi_4 _16591_ (.A1(_07453_),
    .A2(\rbzero.wall_tracer.stepDistY[11] ),
    .B1(_07694_),
    .B2(_09199_),
    .Y(_09200_));
 sky130_fd_sc_hd__nor2_1 _16592_ (.A(_07843_),
    .B(_09200_),
    .Y(_09201_));
 sky130_fd_sc_hd__and2_1 _16593_ (.A(_09052_),
    .B(_09201_),
    .X(_09202_));
 sky130_fd_sc_hd__o22a_1 _16594_ (.A1(_07843_),
    .A2(_09051_),
    .B1(_09200_),
    .B2(_08398_),
    .X(_09203_));
 sky130_fd_sc_hd__nor4_1 _16595_ (.A(_07826_),
    .B(_09197_),
    .C(_09202_),
    .D(_09203_),
    .Y(_09204_));
 sky130_fd_sc_hd__o22a_1 _16596_ (.A1(_07826_),
    .A2(_09197_),
    .B1(_09202_),
    .B2(_09203_),
    .X(_09205_));
 sky130_fd_sc_hd__nor2_1 _16597_ (.A(_09204_),
    .B(_09205_),
    .Y(_09206_));
 sky130_fd_sc_hd__nand2_4 _16598_ (.A(_04938_),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .Y(_09207_));
 sky130_fd_sc_hd__a21oi_1 _16599_ (.A1(_08785_),
    .A2(_09207_),
    .B1(_07835_),
    .Y(_09208_));
 sky130_fd_sc_hd__xnor2_1 _16600_ (.A(_09114_),
    .B(_09208_),
    .Y(_09209_));
 sky130_fd_sc_hd__nor2_1 _16601_ (.A(_07680_),
    .B(_08923_),
    .Y(_09210_));
 sky130_fd_sc_hd__xnor2_1 _16602_ (.A(_09209_),
    .B(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__nand2_1 _16603_ (.A(_09056_),
    .B(_09059_),
    .Y(_09212_));
 sky130_fd_sc_hd__xnor2_1 _16604_ (.A(_09211_),
    .B(_09212_),
    .Y(_09213_));
 sky130_fd_sc_hd__xnor2_1 _16605_ (.A(_09206_),
    .B(_09213_),
    .Y(_09214_));
 sky130_fd_sc_hd__and2_1 _16606_ (.A(_09063_),
    .B(_09065_),
    .X(_09215_));
 sky130_fd_sc_hd__xor2_1 _16607_ (.A(_09214_),
    .B(_09215_),
    .X(_09216_));
 sky130_fd_sc_hd__xnor2_1 _16608_ (.A(_09196_),
    .B(_09216_),
    .Y(_09217_));
 sky130_fd_sc_hd__and2_1 _16609_ (.A(_09069_),
    .B(_09071_),
    .X(_09218_));
 sky130_fd_sc_hd__xor2_1 _16610_ (.A(_09217_),
    .B(_09218_),
    .X(_09219_));
 sky130_fd_sc_hd__xnor2_1 _16611_ (.A(_09181_),
    .B(_09219_),
    .Y(_09220_));
 sky130_fd_sc_hd__and2_1 _16612_ (.A(_09075_),
    .B(_09077_),
    .X(_09221_));
 sky130_fd_sc_hd__xor2_1 _16613_ (.A(_09220_),
    .B(_09221_),
    .X(_09222_));
 sky130_fd_sc_hd__xnor2_1 _16614_ (.A(_09159_),
    .B(_09222_),
    .Y(_09223_));
 sky130_fd_sc_hd__and2_1 _16615_ (.A(_09081_),
    .B(_09083_),
    .X(_09224_));
 sky130_fd_sc_hd__xor2_1 _16616_ (.A(_09223_),
    .B(_09224_),
    .X(_09225_));
 sky130_fd_sc_hd__xnor2_1 _16617_ (.A(_09120_),
    .B(_09225_),
    .Y(_09226_));
 sky130_fd_sc_hd__a21boi_1 _16618_ (.A1(_08974_),
    .A2(_09088_),
    .B1_N(_09087_),
    .Y(_09227_));
 sky130_fd_sc_hd__xor2_1 _16619_ (.A(_09226_),
    .B(_09227_),
    .X(_09228_));
 sky130_fd_sc_hd__xnor2_1 _16620_ (.A(_08972_),
    .B(_09228_),
    .Y(_09229_));
 sky130_fd_sc_hd__and2b_1 _16621_ (.A_N(_09093_),
    .B(_09091_),
    .X(_09230_));
 sky130_fd_sc_hd__a21o_1 _16622_ (.A1(_08844_),
    .A2(_09094_),
    .B1(_09230_),
    .X(_09231_));
 sky130_fd_sc_hd__and2b_1 _16623_ (.A_N(_09229_),
    .B(_09231_),
    .X(_09232_));
 sky130_fd_sc_hd__or2b_1 _16624_ (.A(_09231_),
    .B_N(_09229_),
    .X(_09233_));
 sky130_fd_sc_hd__or2b_2 _16625_ (.A(_09232_),
    .B_N(_09233_),
    .X(_09234_));
 sky130_fd_sc_hd__and2b_1 _16626_ (.A_N(_08955_),
    .B(_09095_),
    .X(_09235_));
 sky130_fd_sc_hd__o21ba_1 _16627_ (.A1(_09096_),
    .A2(_09098_),
    .B1_N(_09235_),
    .X(_09236_));
 sky130_fd_sc_hd__xor2_4 _16628_ (.A(_09234_),
    .B(_09236_),
    .X(_09237_));
 sky130_fd_sc_hd__mux2_1 _16629_ (.A0(\rbzero.debug_overlay.playerY[-1] ),
    .A1(\rbzero.debug_overlay.playerX[-1] ),
    .S(_07343_),
    .X(_09238_));
 sky130_fd_sc_hd__xnor2_1 _16630_ (.A(_08585_),
    .B(_09238_),
    .Y(_09239_));
 sky130_fd_sc_hd__xnor2_1 _16631_ (.A(_09237_),
    .B(_09239_),
    .Y(_09240_));
 sky130_fd_sc_hd__xnor2_1 _16632_ (.A(_09108_),
    .B(_09240_),
    .Y(_09241_));
 sky130_fd_sc_hd__or2_1 _16633_ (.A(\rbzero.wall_tracer.texu[5] ),
    .B(_07338_),
    .X(_09242_));
 sky130_fd_sc_hd__o211a_1 _16634_ (.A1(_04933_),
    .A2(_09241_),
    .B1(_09242_),
    .C1(_07257_),
    .X(_00486_));
 sky130_fd_sc_hd__clkbuf_4 _16635_ (.A(_03292_),
    .X(_09243_));
 sky130_fd_sc_hd__nand2_2 _16636_ (.A(_09243_),
    .B(_03813_),
    .Y(_09244_));
 sky130_fd_sc_hd__nor2_1 _16637_ (.A(_03289_),
    .B(_09244_),
    .Y(_00487_));
 sky130_fd_sc_hd__nor2_4 _16638_ (.A(_03442_),
    .B(_03808_),
    .Y(_09245_));
 sky130_fd_sc_hd__and3_1 _16639_ (.A(_04593_),
    .B(_04087_),
    .C(_09245_),
    .X(_09246_));
 sky130_fd_sc_hd__clkbuf_1 _16640_ (.A(_09246_),
    .X(_00488_));
 sky130_fd_sc_hd__clkbuf_4 _16641_ (.A(_09243_),
    .X(_09247_));
 sky130_fd_sc_hd__or2_1 _16642_ (.A(_04591_),
    .B(_04085_),
    .X(_09248_));
 sky130_fd_sc_hd__and3_1 _16643_ (.A(_09247_),
    .B(_04107_),
    .C(_09248_),
    .X(_09249_));
 sky130_fd_sc_hd__clkbuf_1 _16644_ (.A(_09249_),
    .X(_00489_));
 sky130_fd_sc_hd__nor2_1 _16645_ (.A(_04198_),
    .B(_09244_),
    .Y(_00490_));
 sky130_fd_sc_hd__nor2_1 _16646_ (.A(_04196_),
    .B(_09244_),
    .Y(_00491_));
 sky130_fd_sc_hd__nor2_1 _16647_ (.A(_04220_),
    .B(_09244_),
    .Y(_00492_));
 sky130_fd_sc_hd__nor2_1 _16648_ (.A(_04203_),
    .B(_09244_),
    .Y(_00493_));
 sky130_fd_sc_hd__and3_1 _16649_ (.A(_09247_),
    .B(_03813_),
    .C(_04228_),
    .X(_09250_));
 sky130_fd_sc_hd__clkbuf_1 _16650_ (.A(_09250_),
    .X(_00494_));
 sky130_fd_sc_hd__or2_1 _16651_ (.A(_03294_),
    .B(_04205_),
    .X(_09251_));
 sky130_fd_sc_hd__and3_1 _16652_ (.A(_04206_),
    .B(_09245_),
    .C(_09251_),
    .X(_09252_));
 sky130_fd_sc_hd__clkbuf_1 _16653_ (.A(_09252_),
    .X(_00495_));
 sky130_fd_sc_hd__o21ai_1 _16654_ (.A1(_03296_),
    .A2(_04206_),
    .B1(_09245_),
    .Y(_09253_));
 sky130_fd_sc_hd__a21oi_1 _16655_ (.A1(_03296_),
    .A2(_04206_),
    .B1(_09253_),
    .Y(_00496_));
 sky130_fd_sc_hd__clkbuf_4 _16656_ (.A(_03810_),
    .X(_09254_));
 sky130_fd_sc_hd__buf_2 _16657_ (.A(_09254_),
    .X(_09255_));
 sky130_fd_sc_hd__buf_4 _16658_ (.A(_03728_),
    .X(_09256_));
 sky130_fd_sc_hd__nor2_8 _16659_ (.A(_09256_),
    .B(_03809_),
    .Y(_09257_));
 sky130_fd_sc_hd__clkbuf_4 _16660_ (.A(_09257_),
    .X(_09258_));
 sky130_fd_sc_hd__a22o_1 _16661_ (.A1(\rbzero.row_render.side ),
    .A2(_09255_),
    .B1(_09258_),
    .B2(_07343_),
    .X(_00497_));
 sky130_fd_sc_hd__buf_2 _16662_ (.A(_09257_),
    .X(_09259_));
 sky130_fd_sc_hd__a22o_1 _16663_ (.A1(\rbzero.row_render.size[0] ),
    .A2(_09255_),
    .B1(_07165_),
    .B2(_09259_),
    .X(_00498_));
 sky130_fd_sc_hd__a22o_1 _16664_ (.A1(\rbzero.row_render.size[1] ),
    .A2(_09255_),
    .B1(_07172_),
    .B2(_09259_),
    .X(_00499_));
 sky130_fd_sc_hd__a22o_1 _16665_ (.A1(\rbzero.row_render.size[2] ),
    .A2(_09255_),
    .B1(_07180_),
    .B2(_09259_),
    .X(_00500_));
 sky130_fd_sc_hd__a22o_1 _16666_ (.A1(\rbzero.row_render.size[3] ),
    .A2(_09255_),
    .B1(_07185_),
    .B2(_09259_),
    .X(_00501_));
 sky130_fd_sc_hd__a22o_1 _16667_ (.A1(\rbzero.row_render.size[4] ),
    .A2(_09255_),
    .B1(_07189_),
    .B2(_09259_),
    .X(_00502_));
 sky130_fd_sc_hd__a22o_1 _16668_ (.A1(\rbzero.row_render.size[5] ),
    .A2(_09255_),
    .B1(_07192_),
    .B2(_09259_),
    .X(_00503_));
 sky130_fd_sc_hd__a22o_1 _16669_ (.A1(\rbzero.row_render.size[6] ),
    .A2(_09255_),
    .B1(_07196_),
    .B2(_09259_),
    .X(_00504_));
 sky130_fd_sc_hd__clkbuf_4 _16670_ (.A(_09254_),
    .X(_09260_));
 sky130_fd_sc_hd__a22o_1 _16671_ (.A1(\rbzero.row_render.size[7] ),
    .A2(_09260_),
    .B1(_07199_),
    .B2(_09259_),
    .X(_00505_));
 sky130_fd_sc_hd__a22o_1 _16672_ (.A1(\rbzero.row_render.size[8] ),
    .A2(_09260_),
    .B1(_07202_),
    .B2(_09259_),
    .X(_00506_));
 sky130_fd_sc_hd__a22o_1 _16673_ (.A1(\rbzero.row_render.size[9] ),
    .A2(_09260_),
    .B1(_07206_),
    .B2(_09259_),
    .X(_00507_));
 sky130_fd_sc_hd__buf_4 _16674_ (.A(_09257_),
    .X(_09261_));
 sky130_fd_sc_hd__a22o_1 _16675_ (.A1(\rbzero.row_render.size[10] ),
    .A2(_09260_),
    .B1(_07208_),
    .B2(_09261_),
    .X(_00508_));
 sky130_fd_sc_hd__a22o_1 _16676_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_09260_),
    .B1(_09258_),
    .B2(\rbzero.wall_tracer.texu[0] ),
    .X(_00509_));
 sky130_fd_sc_hd__a22o_1 _16677_ (.A1(\rbzero.row_render.texu[1] ),
    .A2(_09260_),
    .B1(_09258_),
    .B2(\rbzero.wall_tracer.texu[1] ),
    .X(_00510_));
 sky130_fd_sc_hd__a22o_1 _16678_ (.A1(\rbzero.row_render.texu[2] ),
    .A2(_09260_),
    .B1(_09258_),
    .B2(\rbzero.wall_tracer.texu[2] ),
    .X(_00511_));
 sky130_fd_sc_hd__a22o_1 _16679_ (.A1(\rbzero.row_render.texu[3] ),
    .A2(_09260_),
    .B1(_09258_),
    .B2(\rbzero.wall_tracer.texu[3] ),
    .X(_00512_));
 sky130_fd_sc_hd__a22o_1 _16680_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(_09260_),
    .B1(_09258_),
    .B2(\rbzero.wall_tracer.texu[4] ),
    .X(_00513_));
 sky130_fd_sc_hd__a22o_1 _16681_ (.A1(\rbzero.row_render.texu[5] ),
    .A2(_09260_),
    .B1(_09258_),
    .B2(\rbzero.wall_tracer.texu[5] ),
    .X(_00514_));
 sky130_fd_sc_hd__clkbuf_4 _16682_ (.A(_09254_),
    .X(_09262_));
 sky130_fd_sc_hd__a22o_1 _16683_ (.A1(\rbzero.traced_texa[-12] ),
    .A2(_09262_),
    .B1(_09258_),
    .B2(\rbzero.wall_tracer.visualWallDist[-12] ),
    .X(_00515_));
 sky130_fd_sc_hd__a22o_1 _16684_ (.A1(\rbzero.traced_texa[-11] ),
    .A2(_09262_),
    .B1(_09258_),
    .B2(\rbzero.wall_tracer.visualWallDist[-11] ),
    .X(_00516_));
 sky130_fd_sc_hd__buf_2 _16685_ (.A(_09257_),
    .X(_09263_));
 sky130_fd_sc_hd__a22o_1 _16686_ (.A1(\rbzero.traced_texa[-10] ),
    .A2(_09262_),
    .B1(_09263_),
    .B2(\rbzero.wall_tracer.visualWallDist[-10] ),
    .X(_00517_));
 sky130_fd_sc_hd__a22o_1 _16687_ (.A1(\rbzero.traced_texa[-9] ),
    .A2(_09262_),
    .B1(_09263_),
    .B2(\rbzero.wall_tracer.visualWallDist[-9] ),
    .X(_00518_));
 sky130_fd_sc_hd__a22o_1 _16688_ (.A1(\rbzero.traced_texa[-8] ),
    .A2(_09262_),
    .B1(_09263_),
    .B2(\rbzero.wall_tracer.visualWallDist[-8] ),
    .X(_00519_));
 sky130_fd_sc_hd__a22o_1 _16689_ (.A1(\rbzero.traced_texa[-7] ),
    .A2(_09262_),
    .B1(_09263_),
    .B2(\rbzero.wall_tracer.visualWallDist[-7] ),
    .X(_00520_));
 sky130_fd_sc_hd__a22o_1 _16690_ (.A1(\rbzero.traced_texa[-6] ),
    .A2(_09262_),
    .B1(_09263_),
    .B2(\rbzero.wall_tracer.visualWallDist[-6] ),
    .X(_00521_));
 sky130_fd_sc_hd__a22o_1 _16691_ (.A1(\rbzero.traced_texa[-5] ),
    .A2(_09262_),
    .B1(_09263_),
    .B2(\rbzero.wall_tracer.visualWallDist[-5] ),
    .X(_00522_));
 sky130_fd_sc_hd__a22o_1 _16692_ (.A1(\rbzero.traced_texa[-4] ),
    .A2(_09262_),
    .B1(_09263_),
    .B2(\rbzero.wall_tracer.visualWallDist[-4] ),
    .X(_00523_));
 sky130_fd_sc_hd__a22o_1 _16693_ (.A1(\rbzero.traced_texa[-3] ),
    .A2(_09262_),
    .B1(_09263_),
    .B2(\rbzero.wall_tracer.visualWallDist[-3] ),
    .X(_00524_));
 sky130_fd_sc_hd__buf_2 _16694_ (.A(_09254_),
    .X(_09264_));
 sky130_fd_sc_hd__a22o_1 _16695_ (.A1(\rbzero.traced_texa[-2] ),
    .A2(_09264_),
    .B1(_09263_),
    .B2(\rbzero.wall_tracer.visualWallDist[-2] ),
    .X(_00525_));
 sky130_fd_sc_hd__a22o_1 _16696_ (.A1(\rbzero.traced_texa[-1] ),
    .A2(_09264_),
    .B1(_09263_),
    .B2(\rbzero.wall_tracer.visualWallDist[-1] ),
    .X(_00526_));
 sky130_fd_sc_hd__buf_2 _16697_ (.A(_09257_),
    .X(_09265_));
 sky130_fd_sc_hd__a22o_1 _16698_ (.A1(\rbzero.traced_texa[0] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rbzero.wall_tracer.visualWallDist[0] ),
    .X(_00527_));
 sky130_fd_sc_hd__a22o_1 _16699_ (.A1(\rbzero.traced_texa[1] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rbzero.wall_tracer.visualWallDist[1] ),
    .X(_00528_));
 sky130_fd_sc_hd__a22o_1 _16700_ (.A1(\rbzero.traced_texa[2] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rbzero.wall_tracer.visualWallDist[2] ),
    .X(_00529_));
 sky130_fd_sc_hd__a22o_1 _16701_ (.A1(\rbzero.traced_texa[3] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rbzero.wall_tracer.visualWallDist[3] ),
    .X(_00530_));
 sky130_fd_sc_hd__a22o_1 _16702_ (.A1(\rbzero.traced_texa[4] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_00531_));
 sky130_fd_sc_hd__a22o_1 _16703_ (.A1(\rbzero.traced_texa[5] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rbzero.wall_tracer.visualWallDist[5] ),
    .X(_00532_));
 sky130_fd_sc_hd__a22o_1 _16704_ (.A1(\rbzero.traced_texa[6] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rbzero.wall_tracer.visualWallDist[6] ),
    .X(_00533_));
 sky130_fd_sc_hd__a22o_1 _16705_ (.A1(\rbzero.traced_texa[7] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rbzero.wall_tracer.visualWallDist[7] ),
    .X(_00534_));
 sky130_fd_sc_hd__buf_2 _16706_ (.A(_09254_),
    .X(_09266_));
 sky130_fd_sc_hd__a22o_1 _16707_ (.A1(\rbzero.traced_texa[8] ),
    .A2(_09266_),
    .B1(_09265_),
    .B2(\rbzero.wall_tracer.visualWallDist[8] ),
    .X(_00535_));
 sky130_fd_sc_hd__a22o_1 _16708_ (.A1(\rbzero.traced_texa[9] ),
    .A2(_09266_),
    .B1(_09265_),
    .B2(\rbzero.wall_tracer.visualWallDist[9] ),
    .X(_00536_));
 sky130_fd_sc_hd__buf_4 _16709_ (.A(_09257_),
    .X(_09267_));
 sky130_fd_sc_hd__a22o_1 _16710_ (.A1(\rbzero.traced_texa[10] ),
    .A2(_09266_),
    .B1(_09267_),
    .B2(\rbzero.wall_tracer.visualWallDist[10] ),
    .X(_00537_));
 sky130_fd_sc_hd__a22o_1 _16711_ (.A1(\rbzero.traced_texa[11] ),
    .A2(_09266_),
    .B1(_09267_),
    .B2(\rbzero.wall_tracer.visualWallDist[11] ),
    .X(_00538_));
 sky130_fd_sc_hd__or2_1 _16712_ (.A(_03728_),
    .B(_03809_),
    .X(_09268_));
 sky130_fd_sc_hd__clkbuf_4 _16713_ (.A(_09268_),
    .X(_09269_));
 sky130_fd_sc_hd__mux2_1 _16714_ (.A0(\rbzero.wall_tracer.wall[0] ),
    .A1(\rbzero.row_render.wall[0] ),
    .S(_09269_),
    .X(_09270_));
 sky130_fd_sc_hd__clkbuf_1 _16715_ (.A(_09270_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _16716_ (.A0(\rbzero.wall_tracer.wall[1] ),
    .A1(\rbzero.row_render.wall[1] ),
    .S(_09269_),
    .X(_09271_));
 sky130_fd_sc_hd__clkbuf_1 _16717_ (.A(_09271_),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_1 _16718_ (.A0(_04939_),
    .A1(_07254_),
    .S(\rbzero.wall_tracer.state[1] ),
    .X(_09272_));
 sky130_fd_sc_hd__and2_1 _16719_ (.A(_05026_),
    .B(_09272_),
    .X(_09273_));
 sky130_fd_sc_hd__buf_4 _16720_ (.A(_09273_),
    .X(_09274_));
 sky130_fd_sc_hd__clkbuf_4 _16721_ (.A(_09274_),
    .X(_09275_));
 sky130_fd_sc_hd__clkbuf_4 _16722_ (.A(_09275_),
    .X(_09276_));
 sky130_fd_sc_hd__a21oi_1 _16723_ (.A1(_08445_),
    .A2(_08448_),
    .B1(_05121_),
    .Y(_09277_));
 sky130_fd_sc_hd__o21a_1 _16724_ (.A1(_08445_),
    .A2(_08448_),
    .B1(_09277_),
    .X(_09278_));
 sky130_fd_sc_hd__buf_4 _16725_ (.A(_05121_),
    .X(_09279_));
 sky130_fd_sc_hd__nand2_1 _16726_ (.A(\rbzero.wall_tracer.trackDistX[-12] ),
    .B(\rbzero.wall_tracer.stepDistX[-12] ),
    .Y(_09280_));
 sky130_fd_sc_hd__or2_1 _16727_ (.A(\rbzero.wall_tracer.trackDistX[-12] ),
    .B(\rbzero.wall_tracer.stepDistX[-12] ),
    .X(_09281_));
 sky130_fd_sc_hd__nand2_4 _16728_ (.A(_05026_),
    .B(_09272_),
    .Y(_09282_));
 sky130_fd_sc_hd__clkbuf_4 _16729_ (.A(_09282_),
    .X(_09283_));
 sky130_fd_sc_hd__a31o_1 _16730_ (.A1(_09279_),
    .A2(_09280_),
    .A3(_09281_),
    .B1(_09283_),
    .X(_09284_));
 sky130_fd_sc_hd__o22a_1 _16731_ (.A1(\rbzero.wall_tracer.trackDistX[-12] ),
    .A2(_09276_),
    .B1(_09278_),
    .B2(_09284_),
    .X(_00541_));
 sky130_fd_sc_hd__o21a_1 _16732_ (.A1(_08449_),
    .A2(_08322_),
    .B1(_04940_),
    .X(_09285_));
 sky130_fd_sc_hd__a21boi_4 _16733_ (.A1(_08449_),
    .A2(_08322_),
    .B1_N(_09285_),
    .Y(_09286_));
 sky130_fd_sc_hd__or2_1 _16734_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .B(\rbzero.wall_tracer.stepDistX[-11] ),
    .X(_09287_));
 sky130_fd_sc_hd__nand2_1 _16735_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .B(\rbzero.wall_tracer.stepDistX[-11] ),
    .Y(_09288_));
 sky130_fd_sc_hd__nand3b_1 _16736_ (.A_N(_09280_),
    .B(_09287_),
    .C(_09288_),
    .Y(_09289_));
 sky130_fd_sc_hd__a21bo_1 _16737_ (.A1(_09287_),
    .A2(_09288_),
    .B1_N(_09280_),
    .X(_09290_));
 sky130_fd_sc_hd__a31o_1 _16738_ (.A1(_09279_),
    .A2(_09289_),
    .A3(_09290_),
    .B1(_09283_),
    .X(_09291_));
 sky130_fd_sc_hd__o22a_1 _16739_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(_09276_),
    .B1(_09286_),
    .B2(_09291_),
    .X(_00542_));
 sky130_fd_sc_hd__inv_2 _16740_ (.A(_08453_),
    .Y(_09292_));
 sky130_fd_sc_hd__a21oi_1 _16741_ (.A1(_09292_),
    .A2(_08452_),
    .B1(_08450_),
    .Y(_09293_));
 sky130_fd_sc_hd__a211oi_4 _16742_ (.A1(_08450_),
    .A2(_08452_),
    .B1(_09293_),
    .C1(_09279_),
    .Y(_09294_));
 sky130_fd_sc_hd__and2_1 _16743_ (.A(_09288_),
    .B(_09289_),
    .X(_09295_));
 sky130_fd_sc_hd__nor2_1 _16744_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .B(\rbzero.wall_tracer.stepDistX[-10] ),
    .Y(_09296_));
 sky130_fd_sc_hd__and2_1 _16745_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .B(\rbzero.wall_tracer.stepDistX[-10] ),
    .X(_09297_));
 sky130_fd_sc_hd__or3_1 _16746_ (.A(_09295_),
    .B(_09296_),
    .C(_09297_),
    .X(_09298_));
 sky130_fd_sc_hd__o21ai_1 _16747_ (.A1(_09296_),
    .A2(_09297_),
    .B1(_09295_),
    .Y(_09299_));
 sky130_fd_sc_hd__a31o_1 _16748_ (.A1(_09279_),
    .A2(_09298_),
    .A3(_09299_),
    .B1(_09283_),
    .X(_09300_));
 sky130_fd_sc_hd__o22a_1 _16749_ (.A1(\rbzero.wall_tracer.trackDistX[-10] ),
    .A2(_09276_),
    .B1(_09294_),
    .B2(_09300_),
    .X(_00543_));
 sky130_fd_sc_hd__clkbuf_4 _16750_ (.A(_09275_),
    .X(_09301_));
 sky130_fd_sc_hd__and2_1 _16751_ (.A(_07332_),
    .B(_08576_),
    .X(_09302_));
 sky130_fd_sc_hd__buf_4 _16752_ (.A(_05121_),
    .X(_09303_));
 sky130_fd_sc_hd__or2_1 _16753_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .B(\rbzero.wall_tracer.stepDistX[-9] ),
    .X(_09304_));
 sky130_fd_sc_hd__nand2_1 _16754_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .B(\rbzero.wall_tracer.stepDistX[-9] ),
    .Y(_09305_));
 sky130_fd_sc_hd__o21bai_1 _16755_ (.A1(_09295_),
    .A2(_09296_),
    .B1_N(_09297_),
    .Y(_09306_));
 sky130_fd_sc_hd__nand3_1 _16756_ (.A(_09304_),
    .B(_09305_),
    .C(_09306_),
    .Y(_09307_));
 sky130_fd_sc_hd__a21o_1 _16757_ (.A1(_09304_),
    .A2(_09305_),
    .B1(_09306_),
    .X(_09308_));
 sky130_fd_sc_hd__a31o_1 _16758_ (.A1(_09303_),
    .A2(_09307_),
    .A3(_09308_),
    .B1(_09283_),
    .X(_09309_));
 sky130_fd_sc_hd__o22a_1 _16759_ (.A1(\rbzero.wall_tracer.trackDistX[-9] ),
    .A2(_09301_),
    .B1(_09302_),
    .B2(_09309_),
    .X(_00544_));
 sky130_fd_sc_hd__nor2_1 _16760_ (.A(_09279_),
    .B(_08573_),
    .Y(_09310_));
 sky130_fd_sc_hd__nor2_1 _16761_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .Y(_09311_));
 sky130_fd_sc_hd__and2_1 _16762_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .X(_09312_));
 sky130_fd_sc_hd__a21boi_1 _16763_ (.A1(_09304_),
    .A2(_09306_),
    .B1_N(_09305_),
    .Y(_09313_));
 sky130_fd_sc_hd__or3_1 _16764_ (.A(_09311_),
    .B(_09312_),
    .C(_09313_),
    .X(_09314_));
 sky130_fd_sc_hd__o21ai_1 _16765_ (.A1(_09311_),
    .A2(_09312_),
    .B1(_09313_),
    .Y(_09315_));
 sky130_fd_sc_hd__a31o_1 _16766_ (.A1(_09303_),
    .A2(_09314_),
    .A3(_09315_),
    .B1(_09283_),
    .X(_09316_));
 sky130_fd_sc_hd__o22a_1 _16767_ (.A1(\rbzero.wall_tracer.trackDistX[-8] ),
    .A2(_09301_),
    .B1(_09310_),
    .B2(_09316_),
    .X(_00545_));
 sky130_fd_sc_hd__and2_1 _16768_ (.A(_07332_),
    .B(_08571_),
    .X(_09317_));
 sky130_fd_sc_hd__or2_1 _16769_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .X(_09318_));
 sky130_fd_sc_hd__nand2_1 _16770_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .Y(_09319_));
 sky130_fd_sc_hd__o21bai_1 _16771_ (.A1(_09311_),
    .A2(_09313_),
    .B1_N(_09312_),
    .Y(_09320_));
 sky130_fd_sc_hd__nand3_1 _16772_ (.A(_09318_),
    .B(_09319_),
    .C(_09320_),
    .Y(_09321_));
 sky130_fd_sc_hd__a21o_1 _16773_ (.A1(_09318_),
    .A2(_09319_),
    .B1(_09320_),
    .X(_09322_));
 sky130_fd_sc_hd__a31o_1 _16774_ (.A1(_09303_),
    .A2(_09321_),
    .A3(_09322_),
    .B1(_09282_),
    .X(_09323_));
 sky130_fd_sc_hd__o22a_1 _16775_ (.A1(\rbzero.wall_tracer.trackDistX[-7] ),
    .A2(_09301_),
    .B1(_09317_),
    .B2(_09323_),
    .X(_00546_));
 sky130_fd_sc_hd__and2_1 _16776_ (.A(_07332_),
    .B(_08564_),
    .X(_09324_));
 sky130_fd_sc_hd__nor2_1 _16777_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .Y(_09325_));
 sky130_fd_sc_hd__and2_1 _16778_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .X(_09326_));
 sky130_fd_sc_hd__a21boi_1 _16779_ (.A1(_09318_),
    .A2(_09320_),
    .B1_N(_09319_),
    .Y(_09327_));
 sky130_fd_sc_hd__or3_1 _16780_ (.A(_09325_),
    .B(_09326_),
    .C(_09327_),
    .X(_09328_));
 sky130_fd_sc_hd__o21ai_1 _16781_ (.A1(_09325_),
    .A2(_09326_),
    .B1(_09327_),
    .Y(_09329_));
 sky130_fd_sc_hd__a31o_1 _16782_ (.A1(_09303_),
    .A2(_09328_),
    .A3(_09329_),
    .B1(_09282_),
    .X(_09330_));
 sky130_fd_sc_hd__o22a_1 _16783_ (.A1(\rbzero.wall_tracer.trackDistX[-6] ),
    .A2(_09301_),
    .B1(_09324_),
    .B2(_09330_),
    .X(_00547_));
 sky130_fd_sc_hd__nor2_1 _16784_ (.A(_09279_),
    .B(_08700_),
    .Y(_09331_));
 sky130_fd_sc_hd__or2_1 _16785_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .X(_09332_));
 sky130_fd_sc_hd__nand2_1 _16786_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .Y(_09333_));
 sky130_fd_sc_hd__o21bai_1 _16787_ (.A1(_09325_),
    .A2(_09327_),
    .B1_N(_09326_),
    .Y(_09334_));
 sky130_fd_sc_hd__nand3_1 _16788_ (.A(_09332_),
    .B(_09333_),
    .C(_09334_),
    .Y(_09335_));
 sky130_fd_sc_hd__a21o_1 _16789_ (.A1(_09332_),
    .A2(_09333_),
    .B1(_09334_),
    .X(_09336_));
 sky130_fd_sc_hd__a31o_1 _16790_ (.A1(_09303_),
    .A2(_09335_),
    .A3(_09336_),
    .B1(_09282_),
    .X(_09337_));
 sky130_fd_sc_hd__o22a_1 _16791_ (.A1(\rbzero.wall_tracer.trackDistX[-5] ),
    .A2(_09301_),
    .B1(_09331_),
    .B2(_09337_),
    .X(_00548_));
 sky130_fd_sc_hd__nor2_1 _16792_ (.A(_09279_),
    .B(_08828_),
    .Y(_09338_));
 sky130_fd_sc_hd__nor2_1 _16793_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .Y(_09339_));
 sky130_fd_sc_hd__nand2_1 _16794_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .Y(_09340_));
 sky130_fd_sc_hd__and2b_1 _16795_ (.A_N(_09339_),
    .B(_09340_),
    .X(_09341_));
 sky130_fd_sc_hd__a21boi_1 _16796_ (.A1(_09332_),
    .A2(_09334_),
    .B1_N(_09333_),
    .Y(_09342_));
 sky130_fd_sc_hd__xnor2_1 _16797_ (.A(_09341_),
    .B(_09342_),
    .Y(_09343_));
 sky130_fd_sc_hd__a21o_1 _16798_ (.A1(_09279_),
    .A2(_09343_),
    .B1(_09283_),
    .X(_09344_));
 sky130_fd_sc_hd__o22a_1 _16799_ (.A1(\rbzero.wall_tracer.trackDistX[-4] ),
    .A2(_09301_),
    .B1(_09338_),
    .B2(_09344_),
    .X(_00549_));
 sky130_fd_sc_hd__clkbuf_4 _16800_ (.A(_04940_),
    .X(_09345_));
 sky130_fd_sc_hd__or2_1 _16801_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .B(\rbzero.wall_tracer.stepDistX[-3] ),
    .X(_09346_));
 sky130_fd_sc_hd__nand2_1 _16802_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .B(\rbzero.wall_tracer.stepDistX[-3] ),
    .Y(_09347_));
 sky130_fd_sc_hd__o21ai_1 _16803_ (.A1(_09339_),
    .A2(_09342_),
    .B1(_09340_),
    .Y(_09348_));
 sky130_fd_sc_hd__and3_1 _16804_ (.A(_09346_),
    .B(_09347_),
    .C(_09348_),
    .X(_09349_));
 sky130_fd_sc_hd__a21oi_1 _16805_ (.A1(_09346_),
    .A2(_09347_),
    .B1(_09348_),
    .Y(_09350_));
 sky130_fd_sc_hd__clkbuf_4 _16806_ (.A(_04940_),
    .X(_09351_));
 sky130_fd_sc_hd__nand2_1 _16807_ (.A(_09351_),
    .B(_08959_),
    .Y(_09352_));
 sky130_fd_sc_hd__o311a_1 _16808_ (.A1(_09345_),
    .A2(_09349_),
    .A3(_09350_),
    .B1(_09275_),
    .C1(_09352_),
    .X(_09353_));
 sky130_fd_sc_hd__a21oi_1 _16809_ (.A1(_04947_),
    .A2(_09283_),
    .B1(_09353_),
    .Y(_00550_));
 sky130_fd_sc_hd__and2_1 _16810_ (.A(_07332_),
    .B(_09099_),
    .X(_09354_));
 sky130_fd_sc_hd__nor2_1 _16811_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .Y(_09355_));
 sky130_fd_sc_hd__and2_1 _16812_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .X(_09356_));
 sky130_fd_sc_hd__a21boi_1 _16813_ (.A1(_09346_),
    .A2(_09348_),
    .B1_N(_09347_),
    .Y(_09357_));
 sky130_fd_sc_hd__or3_1 _16814_ (.A(_09355_),
    .B(_09356_),
    .C(_09357_),
    .X(_09358_));
 sky130_fd_sc_hd__o21ai_1 _16815_ (.A1(_09355_),
    .A2(_09356_),
    .B1(_09357_),
    .Y(_09359_));
 sky130_fd_sc_hd__a31o_1 _16816_ (.A1(_09303_),
    .A2(_09358_),
    .A3(_09359_),
    .B1(_09282_),
    .X(_09360_));
 sky130_fd_sc_hd__o22a_1 _16817_ (.A1(\rbzero.wall_tracer.trackDistX[-2] ),
    .A2(_09301_),
    .B1(_09354_),
    .B2(_09360_),
    .X(_00551_));
 sky130_fd_sc_hd__nand2_1 _16818_ (.A(_09351_),
    .B(_09237_),
    .Y(_09361_));
 sky130_fd_sc_hd__nor2_1 _16819_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .Y(_09362_));
 sky130_fd_sc_hd__and2_1 _16820_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .X(_09363_));
 sky130_fd_sc_hd__nand2_1 _16821_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .Y(_09364_));
 sky130_fd_sc_hd__o211a_1 _16822_ (.A1(_09362_),
    .A2(_09363_),
    .B1(_09364_),
    .C1(_09358_),
    .X(_09365_));
 sky130_fd_sc_hd__a211oi_2 _16823_ (.A1(_09364_),
    .A2(_09358_),
    .B1(_09362_),
    .C1(_09363_),
    .Y(_09366_));
 sky130_fd_sc_hd__o31a_1 _16824_ (.A1(_07332_),
    .A2(_09365_),
    .A3(_09366_),
    .B1(_09275_),
    .X(_09367_));
 sky130_fd_sc_hd__o2bb2a_1 _16825_ (.A1_N(_09361_),
    .A2_N(_09367_),
    .B1(\rbzero.wall_tracer.trackDistX[-1] ),
    .B2(_09276_),
    .X(_00552_));
 sky130_fd_sc_hd__a21oi_1 _16826_ (.A1(_09235_),
    .A2(_09233_),
    .B1(_09232_),
    .Y(_09368_));
 sky130_fd_sc_hd__o31ai_4 _16827_ (.A1(_09096_),
    .A2(_09098_),
    .A3(_09234_),
    .B1(_09368_),
    .Y(_09369_));
 sky130_fd_sc_hd__or3_1 _16828_ (.A(_09110_),
    .B(_08989_),
    .C(_08990_),
    .X(_09370_));
 sky130_fd_sc_hd__o21ai_1 _16829_ (.A1(_09112_),
    .A2(_09116_),
    .B1(_09370_),
    .Y(_09371_));
 sky130_fd_sc_hd__or2b_1 _16830_ (.A(_09158_),
    .B_N(_09121_),
    .X(_09372_));
 sky130_fd_sc_hd__clkbuf_4 _16831_ (.A(_08979_),
    .X(_09373_));
 sky130_fd_sc_hd__nand2_1 _16832_ (.A(_09124_),
    .B(_09125_),
    .Y(_09374_));
 sky130_fd_sc_hd__o31a_1 _16833_ (.A1(_08429_),
    .A2(_09373_),
    .A3(_09126_),
    .B1(_09374_),
    .X(_09375_));
 sky130_fd_sc_hd__a21oi_2 _16834_ (.A1(_09135_),
    .A2(_09138_),
    .B1(_09375_),
    .Y(_09376_));
 sky130_fd_sc_hd__and3_1 _16835_ (.A(_09135_),
    .B(_09138_),
    .C(_09375_),
    .X(_09377_));
 sky130_fd_sc_hd__or2_1 _16836_ (.A(_09376_),
    .B(_09377_),
    .X(_09378_));
 sky130_fd_sc_hd__a21oi_1 _16837_ (.A1(_09156_),
    .A2(_09372_),
    .B1(_09378_),
    .Y(_09379_));
 sky130_fd_sc_hd__and3_1 _16838_ (.A(_09156_),
    .B(_09372_),
    .C(_09378_),
    .X(_09380_));
 sky130_fd_sc_hd__nor2_1 _16839_ (.A(_09379_),
    .B(_09380_),
    .Y(_09381_));
 sky130_fd_sc_hd__xor2_1 _16840_ (.A(_09371_),
    .B(_09381_),
    .X(_09382_));
 sky130_fd_sc_hd__a21o_1 _16841_ (.A1(_09140_),
    .A2(_09154_),
    .B1(_09152_),
    .X(_09383_));
 sky130_fd_sc_hd__and2b_1 _16842_ (.A_N(_09177_),
    .B(_09162_),
    .X(_09384_));
 sky130_fd_sc_hd__nor2_1 _16843_ (.A(_07878_),
    .B(_08850_),
    .Y(_09385_));
 sky130_fd_sc_hd__nor2_1 _16844_ (.A(_07515_),
    .B(_08978_),
    .Y(_09386_));
 sky130_fd_sc_hd__xnor2_1 _16845_ (.A(_09385_),
    .B(_09386_),
    .Y(_09387_));
 sky130_fd_sc_hd__and3_1 _16846_ (.A(\rbzero.wall_tracer.visualWallDist[11] ),
    .B(_03796_),
    .C(_04929_),
    .X(_09388_));
 sky130_fd_sc_hd__buf_4 _16847_ (.A(_09388_),
    .X(_09389_));
 sky130_fd_sc_hd__nand2_1 _16848_ (.A(_08429_),
    .B(_09389_),
    .Y(_09390_));
 sky130_fd_sc_hd__xor2_1 _16849_ (.A(_09387_),
    .B(_09390_),
    .X(_09391_));
 sky130_fd_sc_hd__or4_1 _16850_ (.A(_08592_),
    .B(_08296_),
    .C(_08716_),
    .D(_08984_),
    .X(_09392_));
 sky130_fd_sc_hd__a2bb2o_1 _16851_ (.A1_N(_08592_),
    .A2_N(_08717_),
    .B1(_08855_),
    .B2(_08507_),
    .X(_09393_));
 sky130_fd_sc_hd__nand2_1 _16852_ (.A(_09392_),
    .B(_09393_),
    .Y(_09394_));
 sky130_fd_sc_hd__nor2_1 _16853_ (.A(_08510_),
    .B(_08722_),
    .Y(_09395_));
 sky130_fd_sc_hd__xor2_1 _16854_ (.A(_09394_),
    .B(_09395_),
    .X(_09396_));
 sky130_fd_sc_hd__o31a_1 _16855_ (.A1(_08510_),
    .A2(_08985_),
    .A3(_09130_),
    .B1(_09131_),
    .X(_09397_));
 sky130_fd_sc_hd__or2_1 _16856_ (.A(_09396_),
    .B(_09397_),
    .X(_09398_));
 sky130_fd_sc_hd__nand2_1 _16857_ (.A(_09396_),
    .B(_09397_),
    .Y(_09399_));
 sky130_fd_sc_hd__and2_1 _16858_ (.A(_09398_),
    .B(_09399_),
    .X(_09400_));
 sky130_fd_sc_hd__nand2_1 _16859_ (.A(_09391_),
    .B(_09400_),
    .Y(_09401_));
 sky130_fd_sc_hd__or2_1 _16860_ (.A(_09391_),
    .B(_09400_),
    .X(_09402_));
 sky130_fd_sc_hd__nand2_1 _16861_ (.A(_09401_),
    .B(_09402_),
    .Y(_09403_));
 sky130_fd_sc_hd__a21bo_1 _16862_ (.A1(_09143_),
    .A2(_09146_),
    .B1_N(_09145_),
    .X(_09404_));
 sky130_fd_sc_hd__or3b_1 _16863_ (.A(_08067_),
    .B(_07685_),
    .C_N(_09028_),
    .X(_09405_));
 sky130_fd_sc_hd__o31a_1 _16864_ (.A1(_08595_),
    .A2(_09166_),
    .A3(_09164_),
    .B1(_09405_),
    .X(_09406_));
 sky130_fd_sc_hd__or4_1 _16865_ (.A(_08086_),
    .B(_08223_),
    .C(_07620_),
    .D(_08671_),
    .X(_09407_));
 sky130_fd_sc_hd__a2bb2o_1 _16866_ (.A1_N(_08086_),
    .A2_N(_07621_),
    .B1(_08536_),
    .B2(_08135_),
    .X(_09408_));
 sky130_fd_sc_hd__nand2_1 _16867_ (.A(_09407_),
    .B(_09408_),
    .Y(_09409_));
 sky130_fd_sc_hd__nor2_1 _16868_ (.A(_08274_),
    .B(_07916_),
    .Y(_09410_));
 sky130_fd_sc_hd__xnor2_1 _16869_ (.A(_09409_),
    .B(_09410_),
    .Y(_09411_));
 sky130_fd_sc_hd__xnor2_1 _16870_ (.A(_09406_),
    .B(_09411_),
    .Y(_09412_));
 sky130_fd_sc_hd__xnor2_1 _16871_ (.A(_09404_),
    .B(_09412_),
    .Y(_09413_));
 sky130_fd_sc_hd__a21oi_1 _16872_ (.A1(_09017_),
    .A2(_09021_),
    .B1(_09147_),
    .Y(_09414_));
 sky130_fd_sc_hd__a21oi_1 _16873_ (.A1(_09141_),
    .A2(_09148_),
    .B1(_09414_),
    .Y(_09415_));
 sky130_fd_sc_hd__nor2_1 _16874_ (.A(_09413_),
    .B(_09415_),
    .Y(_09416_));
 sky130_fd_sc_hd__and2_1 _16875_ (.A(_09413_),
    .B(_09415_),
    .X(_09417_));
 sky130_fd_sc_hd__nor2_1 _16876_ (.A(_09416_),
    .B(_09417_),
    .Y(_09418_));
 sky130_fd_sc_hd__xnor2_1 _16877_ (.A(_09403_),
    .B(_09418_),
    .Y(_09419_));
 sky130_fd_sc_hd__o21ai_1 _16878_ (.A1(_09384_),
    .A2(_09179_),
    .B1(_09419_),
    .Y(_09420_));
 sky130_fd_sc_hd__or3_1 _16879_ (.A(_09384_),
    .B(_09179_),
    .C(_09419_),
    .X(_09421_));
 sky130_fd_sc_hd__nand2_1 _16880_ (.A(_09420_),
    .B(_09421_),
    .Y(_09422_));
 sky130_fd_sc_hd__xnor2_1 _16881_ (.A(_09383_),
    .B(_09422_),
    .Y(_09423_));
 sky130_fd_sc_hd__nor2_1 _16882_ (.A(_09174_),
    .B(_09175_),
    .Y(_09424_));
 sky130_fd_sc_hd__a21o_1 _16883_ (.A1(_09168_),
    .A2(_09176_),
    .B1(_09424_),
    .X(_09425_));
 sky130_fd_sc_hd__or2b_1 _16884_ (.A(_09187_),
    .B_N(_09192_),
    .X(_09426_));
 sky130_fd_sc_hd__or4_1 _16885_ (.A(_07591_),
    .B(_07509_),
    .C(_07685_),
    .D(_07709_),
    .X(_09427_));
 sky130_fd_sc_hd__buf_2 _16886_ (.A(_07509_),
    .X(_09428_));
 sky130_fd_sc_hd__buf_2 _16887_ (.A(_07709_),
    .X(_09429_));
 sky130_fd_sc_hd__a2bb2o_1 _16888_ (.A1_N(_09428_),
    .A2_N(_09429_),
    .B1(_08893_),
    .B2(_09163_),
    .X(_09430_));
 sky130_fd_sc_hd__nand2_1 _16889_ (.A(_09427_),
    .B(_09430_),
    .Y(_09431_));
 sky130_fd_sc_hd__nor2_1 _16890_ (.A(_07598_),
    .B(_09166_),
    .Y(_09432_));
 sky130_fd_sc_hd__xnor2_2 _16891_ (.A(_09431_),
    .B(_09432_),
    .Y(_09433_));
 sky130_fd_sc_hd__and2_1 _16892_ (.A(_07553_),
    .B(_08485_),
    .X(_09434_));
 sky130_fd_sc_hd__nand2_1 _16893_ (.A(_07553_),
    .B(_07837_),
    .Y(_09435_));
 sky130_fd_sc_hd__a22o_1 _16894_ (.A1(_09172_),
    .A2(_09434_),
    .B1(_09435_),
    .B2(_09170_),
    .X(_09436_));
 sky130_fd_sc_hd__or2_1 _16895_ (.A(_07805_),
    .B(_07817_),
    .X(_09437_));
 sky130_fd_sc_hd__xnor2_1 _16896_ (.A(_09436_),
    .B(_09437_),
    .Y(_09438_));
 sky130_fd_sc_hd__or3_1 _16897_ (.A(_07751_),
    .B(_07834_),
    .C(_09170_),
    .X(_09439_));
 sky130_fd_sc_hd__a21boi_1 _16898_ (.A1(_09169_),
    .A2(_09173_),
    .B1_N(_09439_),
    .Y(_09440_));
 sky130_fd_sc_hd__xor2_1 _16899_ (.A(_09438_),
    .B(_09440_),
    .X(_09441_));
 sky130_fd_sc_hd__xnor2_1 _16900_ (.A(_09433_),
    .B(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__a21o_1 _16901_ (.A1(_09426_),
    .A2(_09194_),
    .B1(_09442_),
    .X(_09443_));
 sky130_fd_sc_hd__nand3_1 _16902_ (.A(_09426_),
    .B(_09194_),
    .C(_09442_),
    .Y(_09444_));
 sky130_fd_sc_hd__nand2_1 _16903_ (.A(_09443_),
    .B(_09444_),
    .Y(_09445_));
 sky130_fd_sc_hd__xnor2_1 _16904_ (.A(_09425_),
    .B(_09445_),
    .Y(_09446_));
 sky130_fd_sc_hd__nor2_1 _16905_ (.A(_09047_),
    .B(_09188_),
    .Y(_09447_));
 sky130_fd_sc_hd__a31o_1 _16906_ (.A1(_08771_),
    .A2(_08788_),
    .A3(_09191_),
    .B1(_09447_),
    .X(_09448_));
 sky130_fd_sc_hd__buf_2 _16907_ (.A(_07400_),
    .X(_09449_));
 sky130_fd_sc_hd__and2_1 _16908_ (.A(_08478_),
    .B(_08928_),
    .X(_09450_));
 sky130_fd_sc_hd__buf_2 _16909_ (.A(_09450_),
    .X(_09451_));
 sky130_fd_sc_hd__or3b_1 _16910_ (.A(_09449_),
    .B(_09451_),
    .C_N(_09190_),
    .X(_09452_));
 sky130_fd_sc_hd__o21ai_1 _16911_ (.A1(_09449_),
    .A2(_08917_),
    .B1(_09188_),
    .Y(_09453_));
 sky130_fd_sc_hd__nand2_1 _16912_ (.A(_09452_),
    .B(_09453_),
    .Y(_09454_));
 sky130_fd_sc_hd__nor2_1 _16913_ (.A(_07858_),
    .B(_08780_),
    .Y(_09455_));
 sky130_fd_sc_hd__xnor2_1 _16914_ (.A(_09454_),
    .B(_09455_),
    .Y(_09456_));
 sky130_fd_sc_hd__o21ai_1 _16915_ (.A1(_09202_),
    .A2(_09204_),
    .B1(_09456_),
    .Y(_09457_));
 sky130_fd_sc_hd__or3_1 _16916_ (.A(_09202_),
    .B(_09204_),
    .C(_09456_),
    .X(_09458_));
 sky130_fd_sc_hd__and2_1 _16917_ (.A(_09457_),
    .B(_09458_),
    .X(_09459_));
 sky130_fd_sc_hd__xor2_1 _16918_ (.A(_09448_),
    .B(_09459_),
    .X(_09460_));
 sky130_fd_sc_hd__nand2_1 _16919_ (.A(_08779_),
    .B(_09055_),
    .Y(_09461_));
 sky130_fd_sc_hd__and2_1 _16920_ (.A(_08787_),
    .B(_09207_),
    .X(_09462_));
 sky130_fd_sc_hd__clkbuf_4 _16921_ (.A(_09462_),
    .X(_09463_));
 sky130_fd_sc_hd__or3_1 _16922_ (.A(_07470_),
    .B(_07971_),
    .C(_09200_),
    .X(_09464_));
 sky130_fd_sc_hd__clkbuf_2 _16923_ (.A(_09464_),
    .X(_09465_));
 sky130_fd_sc_hd__o21ai_1 _16924_ (.A1(_08398_),
    .A2(_09200_),
    .B1(_07826_),
    .Y(_09466_));
 sky130_fd_sc_hd__nand2_2 _16925_ (.A(_09465_),
    .B(_09466_),
    .Y(_09467_));
 sky130_fd_sc_hd__nor2_1 _16926_ (.A(_09463_),
    .B(_09467_),
    .Y(_09468_));
 sky130_fd_sc_hd__xnor2_1 _16927_ (.A(_09461_),
    .B(_09468_),
    .Y(_09469_));
 sky130_fd_sc_hd__nand2_4 _16928_ (.A(_04938_),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .Y(_09470_));
 sky130_fd_sc_hd__a21o_1 _16929_ (.A1(_08923_),
    .A2(_09470_),
    .B1(_07835_),
    .X(_09471_));
 sky130_fd_sc_hd__nor2_1 _16930_ (.A(_08335_),
    .B(_09051_),
    .Y(_09472_));
 sky130_fd_sc_hd__xnor2_1 _16931_ (.A(_09471_),
    .B(_09472_),
    .Y(_09473_));
 sky130_fd_sc_hd__or3_1 _16932_ (.A(_07835_),
    .B(_08335_),
    .C(_09200_),
    .X(_09474_));
 sky130_fd_sc_hd__o21ai_1 _16933_ (.A1(_08335_),
    .A2(_09200_),
    .B1(_07835_),
    .Y(_09475_));
 sky130_fd_sc_hd__and3_1 _16934_ (.A(_09201_),
    .B(_09474_),
    .C(_09475_),
    .X(_09476_));
 sky130_fd_sc_hd__o21ba_1 _16935_ (.A1(_09201_),
    .A2(_09473_),
    .B1_N(_09476_),
    .X(_09477_));
 sky130_fd_sc_hd__nand2_1 _16936_ (.A(_09389_),
    .B(_09208_),
    .Y(_09478_));
 sky130_fd_sc_hd__a21boi_1 _16937_ (.A1(_09209_),
    .A2(_09210_),
    .B1_N(_09478_),
    .Y(_09479_));
 sky130_fd_sc_hd__xnor2_1 _16938_ (.A(_09477_),
    .B(_09479_),
    .Y(_09480_));
 sky130_fd_sc_hd__xnor2_1 _16939_ (.A(_09469_),
    .B(_09480_),
    .Y(_09481_));
 sky130_fd_sc_hd__and2b_1 _16940_ (.A_N(_09211_),
    .B(_09212_),
    .X(_09482_));
 sky130_fd_sc_hd__a21o_1 _16941_ (.A1(_09206_),
    .A2(_09213_),
    .B1(_09482_),
    .X(_09483_));
 sky130_fd_sc_hd__xnor2_1 _16942_ (.A(_09481_),
    .B(_09483_),
    .Y(_09484_));
 sky130_fd_sc_hd__xnor2_1 _16943_ (.A(_09460_),
    .B(_09484_),
    .Y(_09485_));
 sky130_fd_sc_hd__nor2_1 _16944_ (.A(_09214_),
    .B(_09215_),
    .Y(_09486_));
 sky130_fd_sc_hd__a21o_1 _16945_ (.A1(_09196_),
    .A2(_09216_),
    .B1(_09486_),
    .X(_09487_));
 sky130_fd_sc_hd__xnor2_1 _16946_ (.A(_09485_),
    .B(_09487_),
    .Y(_09488_));
 sky130_fd_sc_hd__xnor2_1 _16947_ (.A(_09446_),
    .B(_09488_),
    .Y(_09489_));
 sky130_fd_sc_hd__nor2_1 _16948_ (.A(_09217_),
    .B(_09218_),
    .Y(_09490_));
 sky130_fd_sc_hd__a21o_1 _16949_ (.A1(_09181_),
    .A2(_09219_),
    .B1(_09490_),
    .X(_09491_));
 sky130_fd_sc_hd__xnor2_1 _16950_ (.A(_09489_),
    .B(_09491_),
    .Y(_09492_));
 sky130_fd_sc_hd__xnor2_1 _16951_ (.A(_09423_),
    .B(_09492_),
    .Y(_09493_));
 sky130_fd_sc_hd__nor2_1 _16952_ (.A(_09220_),
    .B(_09221_),
    .Y(_09494_));
 sky130_fd_sc_hd__a21oi_1 _16953_ (.A1(_09159_),
    .A2(_09222_),
    .B1(_09494_),
    .Y(_09495_));
 sky130_fd_sc_hd__xor2_1 _16954_ (.A(_09493_),
    .B(_09495_),
    .X(_09496_));
 sky130_fd_sc_hd__xnor2_1 _16955_ (.A(_09382_),
    .B(_09496_),
    .Y(_09497_));
 sky130_fd_sc_hd__nor2_1 _16956_ (.A(_09223_),
    .B(_09224_),
    .Y(_09498_));
 sky130_fd_sc_hd__a21oi_1 _16957_ (.A1(_09120_),
    .A2(_09225_),
    .B1(_09498_),
    .Y(_09499_));
 sky130_fd_sc_hd__xor2_1 _16958_ (.A(_09497_),
    .B(_09499_),
    .X(_09500_));
 sky130_fd_sc_hd__xnor2_1 _16959_ (.A(_09118_),
    .B(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__nor2_1 _16960_ (.A(_09226_),
    .B(_09227_),
    .Y(_09502_));
 sky130_fd_sc_hd__a21oi_1 _16961_ (.A1(_08972_),
    .A2(_09228_),
    .B1(_09502_),
    .Y(_09503_));
 sky130_fd_sc_hd__nor2_1 _16962_ (.A(_09501_),
    .B(_09503_),
    .Y(_09504_));
 sky130_fd_sc_hd__and2_1 _16963_ (.A(_09501_),
    .B(_09503_),
    .X(_09505_));
 sky130_fd_sc_hd__nor2_2 _16964_ (.A(_09504_),
    .B(_09505_),
    .Y(_09506_));
 sky130_fd_sc_hd__xor2_4 _16965_ (.A(_09369_),
    .B(_09506_),
    .X(_09507_));
 sky130_fd_sc_hd__nand2_1 _16966_ (.A(_09351_),
    .B(_09507_),
    .Y(_09508_));
 sky130_fd_sc_hd__or2_1 _16967_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .B(\rbzero.wall_tracer.stepDistX[0] ),
    .X(_09509_));
 sky130_fd_sc_hd__nand2_1 _16968_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .B(\rbzero.wall_tracer.stepDistX[0] ),
    .Y(_09510_));
 sky130_fd_sc_hd__o211a_1 _16969_ (.A1(_09363_),
    .A2(_09366_),
    .B1(_09509_),
    .C1(_09510_),
    .X(_09511_));
 sky130_fd_sc_hd__a211oi_1 _16970_ (.A1(_09509_),
    .A2(_09510_),
    .B1(_09363_),
    .C1(_09366_),
    .Y(_09512_));
 sky130_fd_sc_hd__o31a_1 _16971_ (.A1(_07332_),
    .A2(_09511_),
    .A3(_09512_),
    .B1(_09275_),
    .X(_09513_));
 sky130_fd_sc_hd__o2bb2a_1 _16972_ (.A1_N(_09508_),
    .A2_N(_09513_),
    .B1(\rbzero.wall_tracer.trackDistX[0] ),
    .B2(_09276_),
    .X(_00553_));
 sky130_fd_sc_hd__or2_1 _16973_ (.A(_09497_),
    .B(_09499_),
    .X(_09514_));
 sky130_fd_sc_hd__nand2_1 _16974_ (.A(_09118_),
    .B(_09500_),
    .Y(_09515_));
 sky130_fd_sc_hd__a21o_1 _16975_ (.A1(_09371_),
    .A2(_09381_),
    .B1(_09379_),
    .X(_09516_));
 sky130_fd_sc_hd__or2b_1 _16976_ (.A(_09422_),
    .B_N(_09383_),
    .X(_09517_));
 sky130_fd_sc_hd__nand2_1 _16977_ (.A(_09385_),
    .B(_09386_),
    .Y(_09518_));
 sky130_fd_sc_hd__o21a_1 _16978_ (.A1(_09387_),
    .A2(_09390_),
    .B1(_09518_),
    .X(_09519_));
 sky130_fd_sc_hd__a21oi_2 _16979_ (.A1(_09398_),
    .A2(_09401_),
    .B1(_09519_),
    .Y(_09520_));
 sky130_fd_sc_hd__and3_1 _16980_ (.A(_09398_),
    .B(_09401_),
    .C(_09519_),
    .X(_09521_));
 sky130_fd_sc_hd__or2_1 _16981_ (.A(_09520_),
    .B(_09521_),
    .X(_09522_));
 sky130_fd_sc_hd__a21oi_1 _16982_ (.A1(_09420_),
    .A2(_09517_),
    .B1(_09522_),
    .Y(_09523_));
 sky130_fd_sc_hd__and3_1 _16983_ (.A(_09420_),
    .B(_09517_),
    .C(_09522_),
    .X(_09524_));
 sky130_fd_sc_hd__nor2_1 _16984_ (.A(_09523_),
    .B(_09524_),
    .Y(_09525_));
 sky130_fd_sc_hd__xor2_1 _16985_ (.A(_09376_),
    .B(_09525_),
    .X(_09526_));
 sky130_fd_sc_hd__a31o_1 _16986_ (.A1(_09401_),
    .A2(_09402_),
    .A3(_09418_),
    .B1(_09416_),
    .X(_09527_));
 sky130_fd_sc_hd__or2b_1 _16987_ (.A(_09445_),
    .B_N(_09425_),
    .X(_09528_));
 sky130_fd_sc_hd__or2_1 _16988_ (.A(_07878_),
    .B(_08978_),
    .X(_09529_));
 sky130_fd_sc_hd__nor2_1 _16989_ (.A(_08510_),
    .B(_08850_),
    .Y(_09530_));
 sky130_fd_sc_hd__xnor2_1 _16990_ (.A(_09529_),
    .B(_09530_),
    .Y(_09531_));
 sky130_fd_sc_hd__nor2_1 _16991_ (.A(_07516_),
    .B(_09114_),
    .Y(_09532_));
 sky130_fd_sc_hd__nand2_1 _16992_ (.A(_09531_),
    .B(_09532_),
    .Y(_09533_));
 sky130_fd_sc_hd__or2_1 _16993_ (.A(_09531_),
    .B(_09532_),
    .X(_09534_));
 sky130_fd_sc_hd__and2_1 _16994_ (.A(_09533_),
    .B(_09534_),
    .X(_09535_));
 sky130_fd_sc_hd__o22ai_1 _16995_ (.A1(_08890_),
    .A2(_08718_),
    .B1(_08985_),
    .B2(_08596_),
    .Y(_09536_));
 sky130_fd_sc_hd__or4_1 _16996_ (.A(_08274_),
    .B(_08596_),
    .C(_08718_),
    .D(_08985_),
    .X(_09537_));
 sky130_fd_sc_hd__nand2_1 _16997_ (.A(_09536_),
    .B(_09537_),
    .Y(_09538_));
 sky130_fd_sc_hd__nor2_1 _16998_ (.A(_08599_),
    .B(_08724_),
    .Y(_09539_));
 sky130_fd_sc_hd__xor2_1 _16999_ (.A(_09538_),
    .B(_09539_),
    .X(_09540_));
 sky130_fd_sc_hd__o31a_1 _17000_ (.A1(_08510_),
    .A2(_08724_),
    .A3(_09394_),
    .B1(_09392_),
    .X(_09541_));
 sky130_fd_sc_hd__nor2_1 _17001_ (.A(_09540_),
    .B(_09541_),
    .Y(_09542_));
 sky130_fd_sc_hd__and2_1 _17002_ (.A(_09540_),
    .B(_09541_),
    .X(_09543_));
 sky130_fd_sc_hd__nor2_1 _17003_ (.A(_09542_),
    .B(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__xor2_1 _17004_ (.A(_09535_),
    .B(_09544_),
    .X(_09545_));
 sky130_fd_sc_hd__a21bo_1 _17005_ (.A1(_09408_),
    .A2(_09410_),
    .B1_N(_09407_),
    .X(_09546_));
 sky130_fd_sc_hd__a21bo_1 _17006_ (.A1(_09430_),
    .A2(_09432_),
    .B1_N(_09427_),
    .X(_09547_));
 sky130_fd_sc_hd__or4_1 _17007_ (.A(_08086_),
    .B(_07620_),
    .C(_07936_),
    .D(_08671_),
    .X(_09548_));
 sky130_fd_sc_hd__a2bb2o_1 _17008_ (.A1_N(_07620_),
    .A2_N(_09166_),
    .B1(_08536_),
    .B2(_09018_),
    .X(_09549_));
 sky130_fd_sc_hd__nand2_1 _17009_ (.A(_09548_),
    .B(_09549_),
    .Y(_09550_));
 sky130_fd_sc_hd__nor2_1 _17010_ (.A(_08223_),
    .B(_07916_),
    .Y(_09551_));
 sky130_fd_sc_hd__xnor2_1 _17011_ (.A(_09550_),
    .B(_09551_),
    .Y(_09552_));
 sky130_fd_sc_hd__and2_1 _17012_ (.A(_09547_),
    .B(_09552_),
    .X(_09553_));
 sky130_fd_sc_hd__or2_1 _17013_ (.A(_09547_),
    .B(_09552_),
    .X(_09554_));
 sky130_fd_sc_hd__and2b_1 _17014_ (.A_N(_09553_),
    .B(_09554_),
    .X(_09555_));
 sky130_fd_sc_hd__xnor2_1 _17015_ (.A(_09546_),
    .B(_09555_),
    .Y(_09556_));
 sky130_fd_sc_hd__and2b_1 _17016_ (.A_N(_09406_),
    .B(_09411_),
    .X(_09557_));
 sky130_fd_sc_hd__a21oi_1 _17017_ (.A1(_09404_),
    .A2(_09412_),
    .B1(_09557_),
    .Y(_09558_));
 sky130_fd_sc_hd__nor2_1 _17018_ (.A(_09556_),
    .B(_09558_),
    .Y(_09559_));
 sky130_fd_sc_hd__and2_1 _17019_ (.A(_09556_),
    .B(_09558_),
    .X(_09560_));
 sky130_fd_sc_hd__nor2_1 _17020_ (.A(_09559_),
    .B(_09560_),
    .Y(_09561_));
 sky130_fd_sc_hd__xnor2_1 _17021_ (.A(_09545_),
    .B(_09561_),
    .Y(_09562_));
 sky130_fd_sc_hd__a21oi_1 _17022_ (.A1(_09443_),
    .A2(_09528_),
    .B1(_09562_),
    .Y(_09563_));
 sky130_fd_sc_hd__and3_1 _17023_ (.A(_09443_),
    .B(_09528_),
    .C(_09562_),
    .X(_09564_));
 sky130_fd_sc_hd__nor2_1 _17024_ (.A(_09563_),
    .B(_09564_),
    .Y(_09565_));
 sky130_fd_sc_hd__xor2_1 _17025_ (.A(_09527_),
    .B(_09565_),
    .X(_09566_));
 sky130_fd_sc_hd__nor2_1 _17026_ (.A(_09438_),
    .B(_09440_),
    .Y(_09567_));
 sky130_fd_sc_hd__a21o_1 _17027_ (.A1(_09433_),
    .A2(_09441_),
    .B1(_09567_),
    .X(_09568_));
 sky130_fd_sc_hd__a21bo_1 _17028_ (.A1(_09448_),
    .A2(_09458_),
    .B1_N(_09457_),
    .X(_09569_));
 sky130_fd_sc_hd__or4_1 _17029_ (.A(_07591_),
    .B(_07790_),
    .C(_07672_),
    .D(_07817_),
    .X(_09570_));
 sky130_fd_sc_hd__buf_2 _17030_ (.A(_07672_),
    .X(_09571_));
 sky130_fd_sc_hd__o22ai_1 _17031_ (.A1(_08595_),
    .A2(_09571_),
    .B1(_07817_),
    .B2(_08594_),
    .Y(_09572_));
 sky130_fd_sc_hd__nand2_1 _17032_ (.A(_09570_),
    .B(_09572_),
    .Y(_09573_));
 sky130_fd_sc_hd__nor2_1 _17033_ (.A(_07631_),
    .B(_09429_),
    .Y(_09574_));
 sky130_fd_sc_hd__xnor2_2 _17034_ (.A(_09573_),
    .B(_09574_),
    .Y(_09575_));
 sky130_fd_sc_hd__a21o_1 _17035_ (.A1(_07696_),
    .A2(_08640_),
    .B1(_07800_),
    .X(_09576_));
 sky130_fd_sc_hd__a21oi_2 _17036_ (.A1(_07696_),
    .A2(_08640_),
    .B1(_07890_),
    .Y(_09577_));
 sky130_fd_sc_hd__o22ai_2 _17037_ (.A1(_09170_),
    .A2(_09576_),
    .B1(_09577_),
    .B2(_09434_),
    .Y(_09578_));
 sky130_fd_sc_hd__or2_1 _17038_ (.A(_07805_),
    .B(_07834_),
    .X(_09579_));
 sky130_fd_sc_hd__xnor2_1 _17039_ (.A(_09578_),
    .B(_09579_),
    .Y(_09580_));
 sky130_fd_sc_hd__o2bb2a_1 _17040_ (.A1_N(_09172_),
    .A2_N(_09434_),
    .B1(_09436_),
    .B2(_09437_),
    .X(_09581_));
 sky130_fd_sc_hd__nor2_1 _17041_ (.A(_09580_),
    .B(_09581_),
    .Y(_09582_));
 sky130_fd_sc_hd__nand2_1 _17042_ (.A(_09580_),
    .B(_09581_),
    .Y(_09583_));
 sky130_fd_sc_hd__and2b_1 _17043_ (.A_N(_09582_),
    .B(_09583_),
    .X(_09584_));
 sky130_fd_sc_hd__xor2_1 _17044_ (.A(_09575_),
    .B(_09584_),
    .X(_09585_));
 sky130_fd_sc_hd__and2_1 _17045_ (.A(_09569_),
    .B(_09585_),
    .X(_09586_));
 sky130_fd_sc_hd__or2_1 _17046_ (.A(_09569_),
    .B(_09585_),
    .X(_09587_));
 sky130_fd_sc_hd__or2b_1 _17047_ (.A(_09586_),
    .B_N(_09587_),
    .X(_09588_));
 sky130_fd_sc_hd__xnor2_1 _17048_ (.A(_09568_),
    .B(_09588_),
    .Y(_09589_));
 sky130_fd_sc_hd__o31ai_1 _17049_ (.A1(_09182_),
    .A2(_08780_),
    .A3(_09454_),
    .B1(_09452_),
    .Y(_09590_));
 sky130_fd_sc_hd__o31ai_1 _17050_ (.A1(_09463_),
    .A2(_09461_),
    .A3(_09467_),
    .B1(_09465_),
    .Y(_09591_));
 sky130_fd_sc_hd__or3_1 _17051_ (.A(_09449_),
    .B(_09197_),
    .C(_09188_),
    .X(_09592_));
 sky130_fd_sc_hd__nand2_1 _17052_ (.A(_08046_),
    .B(_09055_),
    .Y(_09593_));
 sky130_fd_sc_hd__o21ai_1 _17053_ (.A1(_09449_),
    .A2(_09451_),
    .B1(_09593_),
    .Y(_09594_));
 sky130_fd_sc_hd__nor2_1 _17054_ (.A(_07858_),
    .B(_08917_),
    .Y(_09595_));
 sky130_fd_sc_hd__nand3_1 _17055_ (.A(_09592_),
    .B(_09594_),
    .C(_09595_),
    .Y(_09596_));
 sky130_fd_sc_hd__a21o_1 _17056_ (.A1(_09592_),
    .A2(_09594_),
    .B1(_09595_),
    .X(_09597_));
 sky130_fd_sc_hd__and3_1 _17057_ (.A(_09591_),
    .B(_09596_),
    .C(_09597_),
    .X(_09598_));
 sky130_fd_sc_hd__a21oi_1 _17058_ (.A1(_09596_),
    .A2(_09597_),
    .B1(_09591_),
    .Y(_09599_));
 sky130_fd_sc_hd__nor2_1 _17059_ (.A(_09598_),
    .B(_09599_),
    .Y(_09600_));
 sky130_fd_sc_hd__xor2_1 _17060_ (.A(_09590_),
    .B(_09600_),
    .X(_09601_));
 sky130_fd_sc_hd__and2_1 _17061_ (.A(_08922_),
    .B(_09470_),
    .X(_09602_));
 sky130_fd_sc_hd__clkbuf_4 _17062_ (.A(_09602_),
    .X(_09603_));
 sky130_fd_sc_hd__or4_1 _17063_ (.A(_07814_),
    .B(_09462_),
    .C(_09467_),
    .D(_09603_),
    .X(_09604_));
 sky130_fd_sc_hd__o22ai_1 _17064_ (.A1(_07814_),
    .A2(_09463_),
    .B1(_09467_),
    .B2(_09603_),
    .Y(_09605_));
 sky130_fd_sc_hd__and2_1 _17065_ (.A(_09604_),
    .B(_09605_),
    .X(_09606_));
 sky130_fd_sc_hd__nand2_1 _17066_ (.A(_08923_),
    .B(_09470_),
    .Y(_09607_));
 sky130_fd_sc_hd__and3_1 _17067_ (.A(_07838_),
    .B(_09607_),
    .C(_09472_),
    .X(_09608_));
 sky130_fd_sc_hd__a21o_1 _17068_ (.A1(_09474_),
    .A2(_09475_),
    .B1(_09201_),
    .X(_09609_));
 sky130_fd_sc_hd__nand2_2 _17069_ (.A(_04939_),
    .B(\rbzero.wall_tracer.stepDistX[10] ),
    .Y(_09610_));
 sky130_fd_sc_hd__o21ai_4 _17070_ (.A1(_04939_),
    .A2(_09051_),
    .B1(_09610_),
    .Y(_09611_));
 sky130_fd_sc_hd__and4b_1 _17071_ (.A_N(_09476_),
    .B(_09608_),
    .C(_09609_),
    .D(_09611_),
    .X(_09612_));
 sky130_fd_sc_hd__a211o_1 _17072_ (.A1(_09609_),
    .A2(_09611_),
    .B1(_09476_),
    .C1(_09608_),
    .X(_09613_));
 sky130_fd_sc_hd__and2b_1 _17073_ (.A_N(_09612_),
    .B(_09613_),
    .X(_09614_));
 sky130_fd_sc_hd__xnor2_1 _17074_ (.A(_09606_),
    .B(_09614_),
    .Y(_09615_));
 sky130_fd_sc_hd__or2b_1 _17075_ (.A(_09479_),
    .B_N(_09477_),
    .X(_09616_));
 sky130_fd_sc_hd__a21bo_1 _17076_ (.A1(_09469_),
    .A2(_09480_),
    .B1_N(_09616_),
    .X(_09617_));
 sky130_fd_sc_hd__xnor2_1 _17077_ (.A(_09615_),
    .B(_09617_),
    .Y(_09618_));
 sky130_fd_sc_hd__xnor2_1 _17078_ (.A(_09601_),
    .B(_09618_),
    .Y(_09619_));
 sky130_fd_sc_hd__or2b_1 _17079_ (.A(_09481_),
    .B_N(_09483_),
    .X(_09620_));
 sky130_fd_sc_hd__a21bo_1 _17080_ (.A1(_09460_),
    .A2(_09484_),
    .B1_N(_09620_),
    .X(_09621_));
 sky130_fd_sc_hd__xnor2_1 _17081_ (.A(_09619_),
    .B(_09621_),
    .Y(_09622_));
 sky130_fd_sc_hd__xnor2_1 _17082_ (.A(_09589_),
    .B(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__or2b_1 _17083_ (.A(_09485_),
    .B_N(_09487_),
    .X(_09624_));
 sky130_fd_sc_hd__a21boi_1 _17084_ (.A1(_09446_),
    .A2(_09488_),
    .B1_N(_09624_),
    .Y(_09625_));
 sky130_fd_sc_hd__xor2_1 _17085_ (.A(_09623_),
    .B(_09625_),
    .X(_09626_));
 sky130_fd_sc_hd__xnor2_1 _17086_ (.A(_09566_),
    .B(_09626_),
    .Y(_09627_));
 sky130_fd_sc_hd__or2b_1 _17087_ (.A(_09489_),
    .B_N(_09491_),
    .X(_09628_));
 sky130_fd_sc_hd__a21boi_1 _17088_ (.A1(_09423_),
    .A2(_09492_),
    .B1_N(_09628_),
    .Y(_09629_));
 sky130_fd_sc_hd__xor2_1 _17089_ (.A(_09627_),
    .B(_09629_),
    .X(_09630_));
 sky130_fd_sc_hd__xnor2_1 _17090_ (.A(_09526_),
    .B(_09630_),
    .Y(_09631_));
 sky130_fd_sc_hd__nor2_1 _17091_ (.A(_09493_),
    .B(_09495_),
    .Y(_09632_));
 sky130_fd_sc_hd__a21oi_1 _17092_ (.A1(_09382_),
    .A2(_09496_),
    .B1(_09632_),
    .Y(_09633_));
 sky130_fd_sc_hd__xnor2_1 _17093_ (.A(_09631_),
    .B(_09633_),
    .Y(_09634_));
 sky130_fd_sc_hd__xor2_1 _17094_ (.A(_09516_),
    .B(_09634_),
    .X(_09635_));
 sky130_fd_sc_hd__and3_1 _17095_ (.A(_09514_),
    .B(_09515_),
    .C(_09635_),
    .X(_09636_));
 sky130_fd_sc_hd__a21o_1 _17096_ (.A1(_09514_),
    .A2(_09515_),
    .B1(_09635_),
    .X(_09637_));
 sky130_fd_sc_hd__and2b_1 _17097_ (.A_N(_09636_),
    .B(_09637_),
    .X(_09638_));
 sky130_fd_sc_hd__a21oi_2 _17098_ (.A1(_09369_),
    .A2(_09506_),
    .B1(_09504_),
    .Y(_09639_));
 sky130_fd_sc_hd__xnor2_4 _17099_ (.A(_09638_),
    .B(_09639_),
    .Y(_09640_));
 sky130_fd_sc_hd__and2_1 _17100_ (.A(_07332_),
    .B(_09640_),
    .X(_09641_));
 sky130_fd_sc_hd__or2_1 _17101_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .B(\rbzero.wall_tracer.stepDistX[1] ),
    .X(_09642_));
 sky130_fd_sc_hd__nand2_1 _17102_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .B(\rbzero.wall_tracer.stepDistX[1] ),
    .Y(_09643_));
 sky130_fd_sc_hd__a21o_1 _17103_ (.A1(\rbzero.wall_tracer.trackDistX[0] ),
    .A2(\rbzero.wall_tracer.stepDistX[0] ),
    .B1(_09511_),
    .X(_09644_));
 sky130_fd_sc_hd__a21o_1 _17104_ (.A1(_09642_),
    .A2(_09643_),
    .B1(_09644_),
    .X(_09645_));
 sky130_fd_sc_hd__and3_1 _17105_ (.A(_09642_),
    .B(_09643_),
    .C(_09644_),
    .X(_09646_));
 sky130_fd_sc_hd__inv_2 _17106_ (.A(_09646_),
    .Y(_09647_));
 sky130_fd_sc_hd__a31o_1 _17107_ (.A1(_09303_),
    .A2(_09645_),
    .A3(_09647_),
    .B1(_09282_),
    .X(_09648_));
 sky130_fd_sc_hd__o22a_1 _17108_ (.A1(\rbzero.wall_tracer.trackDistX[1] ),
    .A2(_09301_),
    .B1(_09641_),
    .B2(_09648_),
    .X(_00554_));
 sky130_fd_sc_hd__or2_1 _17109_ (.A(_09631_),
    .B(_09633_),
    .X(_09649_));
 sky130_fd_sc_hd__or2b_1 _17110_ (.A(_09634_),
    .B_N(_09516_),
    .X(_09650_));
 sky130_fd_sc_hd__a21o_1 _17111_ (.A1(_09376_),
    .A2(_09525_),
    .B1(_09523_),
    .X(_09651_));
 sky130_fd_sc_hd__a21oi_1 _17112_ (.A1(_09527_),
    .A2(_09565_),
    .B1(_09563_),
    .Y(_09652_));
 sky130_fd_sc_hd__a21o_1 _17113_ (.A1(_09535_),
    .A2(_09544_),
    .B1(_09542_),
    .X(_09653_));
 sky130_fd_sc_hd__o31a_1 _17114_ (.A1(_08510_),
    .A2(_08852_),
    .A3(_09529_),
    .B1(_09533_),
    .X(_09654_));
 sky130_fd_sc_hd__inv_2 _17115_ (.A(_09654_),
    .Y(_09655_));
 sky130_fd_sc_hd__nand2_1 _17116_ (.A(_09653_),
    .B(_09655_),
    .Y(_09656_));
 sky130_fd_sc_hd__or2_1 _17117_ (.A(_09653_),
    .B(_09655_),
    .X(_09657_));
 sky130_fd_sc_hd__nand2_1 _17118_ (.A(_09656_),
    .B(_09657_),
    .Y(_09658_));
 sky130_fd_sc_hd__xor2_1 _17119_ (.A(_09652_),
    .B(_09658_),
    .X(_09659_));
 sky130_fd_sc_hd__xor2_1 _17120_ (.A(_09520_),
    .B(_09659_),
    .X(_09660_));
 sky130_fd_sc_hd__a21o_1 _17121_ (.A1(_09545_),
    .A2(_09561_),
    .B1(_09559_),
    .X(_09661_));
 sky130_fd_sc_hd__a21o_1 _17122_ (.A1(_09568_),
    .A2(_09587_),
    .B1(_09586_),
    .X(_09662_));
 sky130_fd_sc_hd__o22ai_1 _17123_ (.A1(_08599_),
    .A2(_08852_),
    .B1(_09373_),
    .B2(_08510_),
    .Y(_09663_));
 sky130_fd_sc_hd__or4_1 _17124_ (.A(_08599_),
    .B(_08510_),
    .C(_08851_),
    .D(_08979_),
    .X(_09664_));
 sky130_fd_sc_hd__nand2_1 _17125_ (.A(_09663_),
    .B(_09664_),
    .Y(_09665_));
 sky130_fd_sc_hd__and3_2 _17126_ (.A(_07505_),
    .B(_07506_),
    .C(_09389_),
    .X(_09666_));
 sky130_fd_sc_hd__xnor2_2 _17127_ (.A(_09665_),
    .B(_09666_),
    .Y(_09667_));
 sky130_fd_sc_hd__a2bb2o_1 _17128_ (.A1_N(_09022_),
    .A2_N(_08718_),
    .B1(_08855_),
    .B2(_08750_),
    .X(_09668_));
 sky130_fd_sc_hd__or4b_1 _17129_ (.A(_09022_),
    .B(_08890_),
    .C(_08718_),
    .D_N(\rbzero.wall_tracer.visualWallDist[7] ),
    .X(_09669_));
 sky130_fd_sc_hd__nand2_1 _17130_ (.A(_09668_),
    .B(_09669_),
    .Y(_09670_));
 sky130_fd_sc_hd__nor2_1 _17131_ (.A(_08596_),
    .B(_08724_),
    .Y(_09671_));
 sky130_fd_sc_hd__xor2_1 _17132_ (.A(_09670_),
    .B(_09671_),
    .X(_09672_));
 sky130_fd_sc_hd__o31a_1 _17133_ (.A1(_08599_),
    .A2(_08725_),
    .A3(_09538_),
    .B1(_09537_),
    .X(_09673_));
 sky130_fd_sc_hd__nor2_1 _17134_ (.A(_09672_),
    .B(_09673_),
    .Y(_09674_));
 sky130_fd_sc_hd__and2_1 _17135_ (.A(_09672_),
    .B(_09673_),
    .X(_09675_));
 sky130_fd_sc_hd__nor2_1 _17136_ (.A(_09674_),
    .B(_09675_),
    .Y(_09676_));
 sky130_fd_sc_hd__xor2_2 _17137_ (.A(_09667_),
    .B(_09676_),
    .X(_09677_));
 sky130_fd_sc_hd__a21bo_1 _17138_ (.A1(_09549_),
    .A2(_09551_),
    .B1_N(_09548_),
    .X(_09678_));
 sky130_fd_sc_hd__a21bo_1 _17139_ (.A1(_09572_),
    .A2(_09574_),
    .B1_N(_09570_),
    .X(_09679_));
 sky130_fd_sc_hd__nor2_1 _17140_ (.A(_07619_),
    .B(_07709_),
    .Y(_09680_));
 sky130_fd_sc_hd__a31o_1 _17141_ (.A1(\rbzero.wall_tracer.visualWallDist[4] ),
    .A2(_03796_),
    .A3(_08123_),
    .B1(_09680_),
    .X(_09681_));
 sky130_fd_sc_hd__or4_1 _17142_ (.A(_07617_),
    .B(_07621_),
    .C(_07709_),
    .D(_09166_),
    .X(_09682_));
 sky130_fd_sc_hd__nand2_1 _17143_ (.A(_09681_),
    .B(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__buf_2 _17144_ (.A(_08086_),
    .X(_09684_));
 sky130_fd_sc_hd__nor2_1 _17145_ (.A(_09684_),
    .B(_08735_),
    .Y(_09685_));
 sky130_fd_sc_hd__xnor2_1 _17146_ (.A(_09683_),
    .B(_09685_),
    .Y(_09686_));
 sky130_fd_sc_hd__and2_1 _17147_ (.A(_09679_),
    .B(_09686_),
    .X(_09687_));
 sky130_fd_sc_hd__or2_1 _17148_ (.A(_09679_),
    .B(_09686_),
    .X(_09688_));
 sky130_fd_sc_hd__and2b_1 _17149_ (.A_N(_09687_),
    .B(_09688_),
    .X(_09689_));
 sky130_fd_sc_hd__xnor2_1 _17150_ (.A(_09678_),
    .B(_09689_),
    .Y(_09690_));
 sky130_fd_sc_hd__a21oi_1 _17151_ (.A1(_09546_),
    .A2(_09555_),
    .B1(_09553_),
    .Y(_09691_));
 sky130_fd_sc_hd__nor2_1 _17152_ (.A(_09690_),
    .B(_09691_),
    .Y(_09692_));
 sky130_fd_sc_hd__and2_1 _17153_ (.A(_09690_),
    .B(_09691_),
    .X(_09693_));
 sky130_fd_sc_hd__nor2_1 _17154_ (.A(_09692_),
    .B(_09693_),
    .Y(_09694_));
 sky130_fd_sc_hd__xor2_2 _17155_ (.A(_09677_),
    .B(_09694_),
    .X(_09695_));
 sky130_fd_sc_hd__xnor2_1 _17156_ (.A(_09662_),
    .B(_09695_),
    .Y(_09696_));
 sky130_fd_sc_hd__xnor2_1 _17157_ (.A(_09661_),
    .B(_09696_),
    .Y(_09697_));
 sky130_fd_sc_hd__a21o_1 _17158_ (.A1(_09575_),
    .A2(_09583_),
    .B1(_09582_),
    .X(_09698_));
 sky130_fd_sc_hd__a21oi_1 _17159_ (.A1(_09590_),
    .A2(_09600_),
    .B1(_09598_),
    .Y(_09699_));
 sky130_fd_sc_hd__nor2_1 _17160_ (.A(_07472_),
    .B(_09428_),
    .Y(_09700_));
 sky130_fd_sc_hd__and3_1 _17161_ (.A(_09163_),
    .B(_07837_),
    .C(_09700_),
    .X(_09701_));
 sky130_fd_sc_hd__a21o_1 _17162_ (.A1(_09163_),
    .A2(_07837_),
    .B1(_09700_),
    .X(_09702_));
 sky130_fd_sc_hd__and2b_1 _17163_ (.A_N(_09701_),
    .B(_09702_),
    .X(_09703_));
 sky130_fd_sc_hd__nor2_1 _17164_ (.A(_07631_),
    .B(_07760_),
    .Y(_09704_));
 sky130_fd_sc_hd__xor2_1 _17165_ (.A(_09703_),
    .B(_09704_),
    .X(_09705_));
 sky130_fd_sc_hd__nor2_1 _17166_ (.A(_08241_),
    .B(_08917_),
    .Y(_09706_));
 sky130_fd_sc_hd__a21o_1 _17167_ (.A1(_07824_),
    .A2(_08793_),
    .B1(_07890_),
    .X(_09707_));
 sky130_fd_sc_hd__a22o_1 _17168_ (.A1(_09577_),
    .A2(_09706_),
    .B1(_09707_),
    .B2(_09576_),
    .X(_09708_));
 sky130_fd_sc_hd__nor2_1 _17169_ (.A(_08760_),
    .B(_08628_),
    .Y(_09709_));
 sky130_fd_sc_hd__xor2_1 _17170_ (.A(_09708_),
    .B(_09709_),
    .X(_09710_));
 sky130_fd_sc_hd__o22a_1 _17171_ (.A1(_09170_),
    .A2(_09576_),
    .B1(_09578_),
    .B2(_09579_),
    .X(_09711_));
 sky130_fd_sc_hd__xor2_1 _17172_ (.A(_09710_),
    .B(_09711_),
    .X(_09712_));
 sky130_fd_sc_hd__nand2_1 _17173_ (.A(_09705_),
    .B(_09712_),
    .Y(_09713_));
 sky130_fd_sc_hd__or2_1 _17174_ (.A(_09705_),
    .B(_09712_),
    .X(_09714_));
 sky130_fd_sc_hd__and2_1 _17175_ (.A(_09713_),
    .B(_09714_),
    .X(_09715_));
 sky130_fd_sc_hd__xnor2_1 _17176_ (.A(_09699_),
    .B(_09715_),
    .Y(_09716_));
 sky130_fd_sc_hd__xor2_1 _17177_ (.A(_09698_),
    .B(_09716_),
    .X(_09717_));
 sky130_fd_sc_hd__nand2_1 _17178_ (.A(_09592_),
    .B(_09596_),
    .Y(_09718_));
 sky130_fd_sc_hd__o41a_1 _17179_ (.A1(_07814_),
    .A2(_09463_),
    .A3(_09467_),
    .A4(_09603_),
    .B1(_09465_),
    .X(_09719_));
 sky130_fd_sc_hd__and2_1 _17180_ (.A(_08771_),
    .B(_09055_),
    .X(_09720_));
 sky130_fd_sc_hd__a21oi_2 _17181_ (.A1(_08787_),
    .A2(_09207_),
    .B1(_08272_),
    .Y(_09721_));
 sky130_fd_sc_hd__a21o_1 _17182_ (.A1(_08787_),
    .A2(_09207_),
    .B1(_09449_),
    .X(_09722_));
 sky130_fd_sc_hd__o22a_1 _17183_ (.A1(_09720_),
    .A2(_09721_),
    .B1(_09722_),
    .B2(_09593_),
    .X(_09723_));
 sky130_fd_sc_hd__nor2_1 _17184_ (.A(_07858_),
    .B(_09451_),
    .Y(_09724_));
 sky130_fd_sc_hd__xor2_1 _17185_ (.A(_09723_),
    .B(_09724_),
    .X(_09725_));
 sky130_fd_sc_hd__xnor2_1 _17186_ (.A(_09719_),
    .B(_09725_),
    .Y(_09726_));
 sky130_fd_sc_hd__xor2_1 _17187_ (.A(_09718_),
    .B(_09726_),
    .X(_09727_));
 sky130_fd_sc_hd__nand2_1 _17188_ (.A(_08779_),
    .B(_09611_),
    .Y(_09728_));
 sky130_fd_sc_hd__a32o_1 _17189_ (.A1(_09465_),
    .A2(_09466_),
    .A3(_09611_),
    .B1(_09607_),
    .B2(_08779_),
    .X(_09729_));
 sky130_fd_sc_hd__o31a_1 _17190_ (.A1(_09467_),
    .A2(_09603_),
    .A3(_09728_),
    .B1(_09729_),
    .X(_09730_));
 sky130_fd_sc_hd__nand2_2 _17191_ (.A(_04938_),
    .B(\rbzero.wall_tracer.stepDistX[11] ),
    .Y(_09731_));
 sky130_fd_sc_hd__o21ai_2 _17192_ (.A1(_04939_),
    .A2(_09200_),
    .B1(_09731_),
    .Y(_09732_));
 sky130_fd_sc_hd__or4bb_2 _17193_ (.A(_09474_),
    .B(_09476_),
    .C_N(_09609_),
    .D_N(_09732_),
    .X(_09733_));
 sky130_fd_sc_hd__inv_2 _17194_ (.A(_09474_),
    .Y(_09734_));
 sky130_fd_sc_hd__a211o_2 _17195_ (.A1(_09609_),
    .A2(_09732_),
    .B1(_09734_),
    .C1(_09476_),
    .X(_09735_));
 sky130_fd_sc_hd__nand2_1 _17196_ (.A(_09733_),
    .B(_09735_),
    .Y(_09736_));
 sky130_fd_sc_hd__xor2_1 _17197_ (.A(_09730_),
    .B(_09736_),
    .X(_09737_));
 sky130_fd_sc_hd__a21oi_1 _17198_ (.A1(_09606_),
    .A2(_09613_),
    .B1(_09612_),
    .Y(_09738_));
 sky130_fd_sc_hd__xor2_1 _17199_ (.A(_09737_),
    .B(_09738_),
    .X(_09739_));
 sky130_fd_sc_hd__xnor2_1 _17200_ (.A(_09727_),
    .B(_09739_),
    .Y(_09740_));
 sky130_fd_sc_hd__or2b_1 _17201_ (.A(_09615_),
    .B_N(_09617_),
    .X(_09741_));
 sky130_fd_sc_hd__a21bo_1 _17202_ (.A1(_09601_),
    .A2(_09618_),
    .B1_N(_09741_),
    .X(_09742_));
 sky130_fd_sc_hd__xnor2_1 _17203_ (.A(_09740_),
    .B(_09742_),
    .Y(_09743_));
 sky130_fd_sc_hd__xnor2_1 _17204_ (.A(_09717_),
    .B(_09743_),
    .Y(_09744_));
 sky130_fd_sc_hd__or2b_1 _17205_ (.A(_09619_),
    .B_N(_09621_),
    .X(_09745_));
 sky130_fd_sc_hd__a21boi_1 _17206_ (.A1(_09589_),
    .A2(_09622_),
    .B1_N(_09745_),
    .Y(_09746_));
 sky130_fd_sc_hd__xor2_1 _17207_ (.A(_09744_),
    .B(_09746_),
    .X(_09747_));
 sky130_fd_sc_hd__xnor2_1 _17208_ (.A(_09697_),
    .B(_09747_),
    .Y(_09748_));
 sky130_fd_sc_hd__nor2_1 _17209_ (.A(_09623_),
    .B(_09625_),
    .Y(_09749_));
 sky130_fd_sc_hd__a21oi_1 _17210_ (.A1(_09566_),
    .A2(_09626_),
    .B1(_09749_),
    .Y(_09750_));
 sky130_fd_sc_hd__xor2_1 _17211_ (.A(_09748_),
    .B(_09750_),
    .X(_09751_));
 sky130_fd_sc_hd__xnor2_1 _17212_ (.A(_09660_),
    .B(_09751_),
    .Y(_09752_));
 sky130_fd_sc_hd__nor2_1 _17213_ (.A(_09627_),
    .B(_09629_),
    .Y(_09753_));
 sky130_fd_sc_hd__a21oi_1 _17214_ (.A1(_09526_),
    .A2(_09630_),
    .B1(_09753_),
    .Y(_09754_));
 sky130_fd_sc_hd__xor2_1 _17215_ (.A(_09752_),
    .B(_09754_),
    .X(_09755_));
 sky130_fd_sc_hd__xnor2_1 _17216_ (.A(_09651_),
    .B(_09755_),
    .Y(_09756_));
 sky130_fd_sc_hd__a21o_1 _17217_ (.A1(_09649_),
    .A2(_09650_),
    .B1(_09756_),
    .X(_09757_));
 sky130_fd_sc_hd__and3_1 _17218_ (.A(_09649_),
    .B(_09650_),
    .C(_09756_),
    .X(_09758_));
 sky130_fd_sc_hd__inv_2 _17219_ (.A(_09758_),
    .Y(_09759_));
 sky130_fd_sc_hd__nand2_2 _17220_ (.A(_09757_),
    .B(_09759_),
    .Y(_09760_));
 sky130_fd_sc_hd__and2_1 _17221_ (.A(_09506_),
    .B(_09638_),
    .X(_09761_));
 sky130_fd_sc_hd__o31a_1 _17222_ (.A1(_09501_),
    .A2(_09503_),
    .A3(_09636_),
    .B1(_09637_),
    .X(_09762_));
 sky130_fd_sc_hd__a21bo_1 _17223_ (.A1(_09369_),
    .A2(_09761_),
    .B1_N(_09762_),
    .X(_09763_));
 sky130_fd_sc_hd__xnor2_4 _17224_ (.A(_09760_),
    .B(_09763_),
    .Y(_09764_));
 sky130_fd_sc_hd__and2_1 _17225_ (.A(_09345_),
    .B(_09764_),
    .X(_09765_));
 sky130_fd_sc_hd__nand2_1 _17226_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .B(\rbzero.wall_tracer.stepDistX[2] ),
    .Y(_09766_));
 sky130_fd_sc_hd__or2_1 _17227_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .B(\rbzero.wall_tracer.stepDistX[2] ),
    .X(_09767_));
 sky130_fd_sc_hd__nand2_1 _17228_ (.A(_09643_),
    .B(_09647_),
    .Y(_09768_));
 sky130_fd_sc_hd__and3_1 _17229_ (.A(_09766_),
    .B(_09767_),
    .C(_09768_),
    .X(_09769_));
 sky130_fd_sc_hd__inv_2 _17230_ (.A(_09769_),
    .Y(_09770_));
 sky130_fd_sc_hd__a21o_1 _17231_ (.A1(_09766_),
    .A2(_09767_),
    .B1(_09768_),
    .X(_09771_));
 sky130_fd_sc_hd__a31o_1 _17232_ (.A1(_09303_),
    .A2(_09770_),
    .A3(_09771_),
    .B1(_09282_),
    .X(_09772_));
 sky130_fd_sc_hd__o22a_1 _17233_ (.A1(\rbzero.wall_tracer.trackDistX[2] ),
    .A2(_09301_),
    .B1(_09765_),
    .B2(_09772_),
    .X(_00555_));
 sky130_fd_sc_hd__or2_1 _17234_ (.A(_09752_),
    .B(_09754_),
    .X(_09773_));
 sky130_fd_sc_hd__nand2_1 _17235_ (.A(_09651_),
    .B(_09755_),
    .Y(_09774_));
 sky130_fd_sc_hd__nand2_1 _17236_ (.A(_09520_),
    .B(_09659_),
    .Y(_09775_));
 sky130_fd_sc_hd__o21ai_1 _17237_ (.A1(_09652_),
    .A2(_09658_),
    .B1(_09775_),
    .Y(_09776_));
 sky130_fd_sc_hd__nand2_1 _17238_ (.A(_09662_),
    .B(_09695_),
    .Y(_09777_));
 sky130_fd_sc_hd__or2b_1 _17239_ (.A(_09696_),
    .B_N(_09661_),
    .X(_09778_));
 sky130_fd_sc_hd__a21o_1 _17240_ (.A1(_09667_),
    .A2(_09676_),
    .B1(_09674_),
    .X(_09779_));
 sky130_fd_sc_hd__a21boi_1 _17241_ (.A1(_09663_),
    .A2(_09666_),
    .B1_N(_09664_),
    .Y(_09780_));
 sky130_fd_sc_hd__inv_2 _17242_ (.A(_09780_),
    .Y(_09781_));
 sky130_fd_sc_hd__nand2_1 _17243_ (.A(_09779_),
    .B(_09781_),
    .Y(_09782_));
 sky130_fd_sc_hd__or2_1 _17244_ (.A(_09779_),
    .B(_09781_),
    .X(_09783_));
 sky130_fd_sc_hd__nand2_1 _17245_ (.A(_09782_),
    .B(_09783_),
    .Y(_09784_));
 sky130_fd_sc_hd__a21oi_1 _17246_ (.A1(_09777_),
    .A2(_09778_),
    .B1(_09784_),
    .Y(_09785_));
 sky130_fd_sc_hd__and3_1 _17247_ (.A(_09777_),
    .B(_09778_),
    .C(_09784_),
    .X(_09786_));
 sky130_fd_sc_hd__nor2_1 _17248_ (.A(_09785_),
    .B(_09786_),
    .Y(_09787_));
 sky130_fd_sc_hd__xnor2_1 _17249_ (.A(_09656_),
    .B(_09787_),
    .Y(_09788_));
 sky130_fd_sc_hd__a21o_1 _17250_ (.A1(_09677_),
    .A2(_09694_),
    .B1(_09692_),
    .X(_09789_));
 sky130_fd_sc_hd__or2b_1 _17251_ (.A(_09699_),
    .B_N(_09715_),
    .X(_09790_));
 sky130_fd_sc_hd__a21bo_1 _17252_ (.A1(_09698_),
    .A2(_09716_),
    .B1_N(_09790_),
    .X(_09791_));
 sky130_fd_sc_hd__o22a_1 _17253_ (.A1(_08596_),
    .A2(_08851_),
    .B1(_09373_),
    .B2(_08599_),
    .X(_09792_));
 sky130_fd_sc_hd__or4_1 _17254_ (.A(_08596_),
    .B(_08599_),
    .C(_08851_),
    .D(_08979_),
    .X(_09793_));
 sky130_fd_sc_hd__or2b_1 _17255_ (.A(_09792_),
    .B_N(_09793_),
    .X(_09794_));
 sky130_fd_sc_hd__nor2_1 _17256_ (.A(_07882_),
    .B(_09115_),
    .Y(_09795_));
 sky130_fd_sc_hd__xnor2_1 _17257_ (.A(_09794_),
    .B(_09795_),
    .Y(_09796_));
 sky130_fd_sc_hd__nor2_1 _17258_ (.A(_09684_),
    .B(_08717_),
    .Y(_09797_));
 sky130_fd_sc_hd__a21oi_1 _17259_ (.A1(_08135_),
    .A2(_08855_),
    .B1(_09797_),
    .Y(_09798_));
 sky130_fd_sc_hd__or4_1 _17260_ (.A(_09684_),
    .B(_09022_),
    .C(_08718_),
    .D(_08985_),
    .X(_09799_));
 sky130_fd_sc_hd__or2b_1 _17261_ (.A(_09798_),
    .B_N(_09799_),
    .X(_09800_));
 sky130_fd_sc_hd__nor2_1 _17262_ (.A(_08890_),
    .B(_08725_),
    .Y(_09801_));
 sky130_fd_sc_hd__xor2_1 _17263_ (.A(_09800_),
    .B(_09801_),
    .X(_09802_));
 sky130_fd_sc_hd__o31a_1 _17264_ (.A1(_08596_),
    .A2(_08725_),
    .A3(_09670_),
    .B1(_09669_),
    .X(_09803_));
 sky130_fd_sc_hd__nor2_1 _17265_ (.A(_09802_),
    .B(_09803_),
    .Y(_09804_));
 sky130_fd_sc_hd__and2_1 _17266_ (.A(_09802_),
    .B(_09803_),
    .X(_09805_));
 sky130_fd_sc_hd__nor2_1 _17267_ (.A(_09804_),
    .B(_09805_),
    .Y(_09806_));
 sky130_fd_sc_hd__xor2_1 _17268_ (.A(_09796_),
    .B(_09806_),
    .X(_09807_));
 sky130_fd_sc_hd__a21bo_1 _17269_ (.A1(_09681_),
    .A2(_09685_),
    .B1_N(_09682_),
    .X(_09808_));
 sky130_fd_sc_hd__a21oi_1 _17270_ (.A1(_09702_),
    .A2(_09704_),
    .B1(_09701_),
    .Y(_09809_));
 sky130_fd_sc_hd__or4_1 _17271_ (.A(_07618_),
    .B(_08732_),
    .C(_09571_),
    .D(_09429_),
    .X(_09810_));
 sky130_fd_sc_hd__o22ai_1 _17272_ (.A1(_08732_),
    .A2(_09571_),
    .B1(_09429_),
    .B2(_07618_),
    .Y(_09811_));
 sky130_fd_sc_hd__nand2_1 _17273_ (.A(_09810_),
    .B(_09811_),
    .Y(_09812_));
 sky130_fd_sc_hd__nor2_1 _17274_ (.A(_09166_),
    .B(_08735_),
    .Y(_09813_));
 sky130_fd_sc_hd__xor2_1 _17275_ (.A(_09812_),
    .B(_09813_),
    .X(_09814_));
 sky130_fd_sc_hd__nor2_1 _17276_ (.A(_09809_),
    .B(_09814_),
    .Y(_09815_));
 sky130_fd_sc_hd__nand2_1 _17277_ (.A(_09809_),
    .B(_09814_),
    .Y(_09816_));
 sky130_fd_sc_hd__and2b_1 _17278_ (.A_N(_09815_),
    .B(_09816_),
    .X(_09817_));
 sky130_fd_sc_hd__xnor2_1 _17279_ (.A(_09808_),
    .B(_09817_),
    .Y(_09818_));
 sky130_fd_sc_hd__a21oi_1 _17280_ (.A1(_09678_),
    .A2(_09689_),
    .B1(_09687_),
    .Y(_09819_));
 sky130_fd_sc_hd__nor2_1 _17281_ (.A(_09818_),
    .B(_09819_),
    .Y(_09820_));
 sky130_fd_sc_hd__and2_1 _17282_ (.A(_09818_),
    .B(_09819_),
    .X(_09821_));
 sky130_fd_sc_hd__nor2_1 _17283_ (.A(_09820_),
    .B(_09821_),
    .Y(_09822_));
 sky130_fd_sc_hd__xor2_1 _17284_ (.A(_09807_),
    .B(_09822_),
    .X(_09823_));
 sky130_fd_sc_hd__xnor2_1 _17285_ (.A(_09791_),
    .B(_09823_),
    .Y(_09824_));
 sky130_fd_sc_hd__xnor2_1 _17286_ (.A(_09789_),
    .B(_09824_),
    .Y(_09825_));
 sky130_fd_sc_hd__o21ai_1 _17287_ (.A1(_09710_),
    .A2(_09711_),
    .B1(_09713_),
    .Y(_09826_));
 sky130_fd_sc_hd__and2b_1 _17288_ (.A_N(_09719_),
    .B(_09725_),
    .X(_09827_));
 sky130_fd_sc_hd__a21oi_1 _17289_ (.A1(_09718_),
    .A2(_09726_),
    .B1(_09827_),
    .Y(_09828_));
 sky130_fd_sc_hd__a21oi_4 _17290_ (.A1(_04933_),
    .A2(_07648_),
    .B1(_07650_),
    .Y(_09829_));
 sky130_fd_sc_hd__or4_1 _17291_ (.A(_08594_),
    .B(_08595_),
    .C(_09829_),
    .D(_08628_),
    .X(_09830_));
 sky130_fd_sc_hd__a22o_1 _17292_ (.A1(_07520_),
    .A2(_07651_),
    .B1(_08636_),
    .B2(_09163_),
    .X(_09831_));
 sky130_fd_sc_hd__nand2_1 _17293_ (.A(_09830_),
    .B(_09831_),
    .Y(_09832_));
 sky130_fd_sc_hd__buf_2 _17294_ (.A(_07472_),
    .X(_09833_));
 sky130_fd_sc_hd__nor2_1 _17295_ (.A(_09833_),
    .B(_07631_),
    .Y(_09834_));
 sky130_fd_sc_hd__xnor2_1 _17296_ (.A(_09832_),
    .B(_09834_),
    .Y(_09835_));
 sky130_fd_sc_hd__nor2_1 _17297_ (.A(_08240_),
    .B(_09451_),
    .Y(_09836_));
 sky130_fd_sc_hd__or3_1 _17298_ (.A(_07800_),
    .B(_09451_),
    .C(_09707_),
    .X(_09837_));
 sky130_fd_sc_hd__o21ai_1 _17299_ (.A1(_09706_),
    .A2(_09836_),
    .B1(_09837_),
    .Y(_09838_));
 sky130_fd_sc_hd__nor2_1 _17300_ (.A(_08760_),
    .B(_08780_),
    .Y(_09839_));
 sky130_fd_sc_hd__xor2_1 _17301_ (.A(_09838_),
    .B(_09839_),
    .X(_09840_));
 sky130_fd_sc_hd__nand2_1 _17302_ (.A(_09577_),
    .B(_09706_),
    .Y(_09841_));
 sky130_fd_sc_hd__o31a_1 _17303_ (.A1(_08760_),
    .A2(_08628_),
    .A3(_09708_),
    .B1(_09841_),
    .X(_09842_));
 sky130_fd_sc_hd__xor2_1 _17304_ (.A(_09840_),
    .B(_09842_),
    .X(_09843_));
 sky130_fd_sc_hd__xnor2_1 _17305_ (.A(_09835_),
    .B(_09843_),
    .Y(_09844_));
 sky130_fd_sc_hd__xor2_1 _17306_ (.A(_09828_),
    .B(_09844_),
    .X(_09845_));
 sky130_fd_sc_hd__nand2_1 _17307_ (.A(_09826_),
    .B(_09845_),
    .Y(_09846_));
 sky130_fd_sc_hd__or2_1 _17308_ (.A(_09826_),
    .B(_09845_),
    .X(_09847_));
 sky130_fd_sc_hd__and2_1 _17309_ (.A(_09846_),
    .B(_09847_),
    .X(_09848_));
 sky130_fd_sc_hd__a2bb2o_1 _17310_ (.A1_N(_09593_),
    .A2_N(_09722_),
    .B1(_09723_),
    .B2(_09724_),
    .X(_09849_));
 sky130_fd_sc_hd__o31a_1 _17311_ (.A1(_09467_),
    .A2(_09603_),
    .A3(_09728_),
    .B1(_09465_),
    .X(_09850_));
 sky130_fd_sc_hd__a21o_1 _17312_ (.A1(_08923_),
    .A2(_09470_),
    .B1(_08272_),
    .X(_09851_));
 sky130_fd_sc_hd__a32oi_2 _17313_ (.A1(_08771_),
    .A2(_09607_),
    .A3(_09721_),
    .B1(_09722_),
    .B2(_09851_),
    .Y(_09852_));
 sky130_fd_sc_hd__nor2_1 _17314_ (.A(_09182_),
    .B(_09197_),
    .Y(_09853_));
 sky130_fd_sc_hd__xnor2_1 _17315_ (.A(_09852_),
    .B(_09853_),
    .Y(_09854_));
 sky130_fd_sc_hd__xor2_1 _17316_ (.A(_09850_),
    .B(_09854_),
    .X(_09855_));
 sky130_fd_sc_hd__xor2_1 _17317_ (.A(_09849_),
    .B(_09855_),
    .X(_09856_));
 sky130_fd_sc_hd__and3_1 _17318_ (.A(_09465_),
    .B(_09466_),
    .C(_09732_),
    .X(_09857_));
 sky130_fd_sc_hd__xnor2_1 _17319_ (.A(_09728_),
    .B(_09857_),
    .Y(_09858_));
 sky130_fd_sc_hd__nand3_1 _17320_ (.A(_09733_),
    .B(_09735_),
    .C(_09858_),
    .Y(_09859_));
 sky130_fd_sc_hd__a21o_1 _17321_ (.A1(_09733_),
    .A2(_09735_),
    .B1(_09858_),
    .X(_09860_));
 sky130_fd_sc_hd__and4b_2 _17322_ (.A_N(_09476_),
    .B(_09609_),
    .C(_09732_),
    .D(_09734_),
    .X(_09861_));
 sky130_fd_sc_hd__a21o_1 _17323_ (.A1(_09730_),
    .A2(_09735_),
    .B1(_09861_),
    .X(_09862_));
 sky130_fd_sc_hd__and3_1 _17324_ (.A(_09859_),
    .B(_09860_),
    .C(_09862_),
    .X(_09863_));
 sky130_fd_sc_hd__a21o_1 _17325_ (.A1(_09859_),
    .A2(_09860_),
    .B1(_09862_),
    .X(_09864_));
 sky130_fd_sc_hd__and2b_1 _17326_ (.A_N(_09863_),
    .B(_09864_),
    .X(_09865_));
 sky130_fd_sc_hd__xor2_1 _17327_ (.A(_09856_),
    .B(_09865_),
    .X(_09866_));
 sky130_fd_sc_hd__nor2_1 _17328_ (.A(_09737_),
    .B(_09738_),
    .Y(_09867_));
 sky130_fd_sc_hd__a21o_1 _17329_ (.A1(_09727_),
    .A2(_09739_),
    .B1(_09867_),
    .X(_09868_));
 sky130_fd_sc_hd__xor2_1 _17330_ (.A(_09866_),
    .B(_09868_),
    .X(_09869_));
 sky130_fd_sc_hd__xnor2_1 _17331_ (.A(_09848_),
    .B(_09869_),
    .Y(_09870_));
 sky130_fd_sc_hd__or2b_1 _17332_ (.A(_09740_),
    .B_N(_09742_),
    .X(_09871_));
 sky130_fd_sc_hd__a21boi_1 _17333_ (.A1(_09717_),
    .A2(_09743_),
    .B1_N(_09871_),
    .Y(_09872_));
 sky130_fd_sc_hd__xor2_1 _17334_ (.A(_09870_),
    .B(_09872_),
    .X(_09873_));
 sky130_fd_sc_hd__xnor2_1 _17335_ (.A(_09825_),
    .B(_09873_),
    .Y(_09874_));
 sky130_fd_sc_hd__nor2_1 _17336_ (.A(_09744_),
    .B(_09746_),
    .Y(_09875_));
 sky130_fd_sc_hd__a21oi_1 _17337_ (.A1(_09697_),
    .A2(_09747_),
    .B1(_09875_),
    .Y(_09876_));
 sky130_fd_sc_hd__xor2_1 _17338_ (.A(_09874_),
    .B(_09876_),
    .X(_09877_));
 sky130_fd_sc_hd__xnor2_1 _17339_ (.A(_09788_),
    .B(_09877_),
    .Y(_09878_));
 sky130_fd_sc_hd__nor2_1 _17340_ (.A(_09748_),
    .B(_09750_),
    .Y(_09879_));
 sky130_fd_sc_hd__a21oi_1 _17341_ (.A1(_09660_),
    .A2(_09751_),
    .B1(_09879_),
    .Y(_09880_));
 sky130_fd_sc_hd__xnor2_1 _17342_ (.A(_09878_),
    .B(_09880_),
    .Y(_09881_));
 sky130_fd_sc_hd__xor2_1 _17343_ (.A(_09776_),
    .B(_09881_),
    .X(_09882_));
 sky130_fd_sc_hd__and3_1 _17344_ (.A(_09773_),
    .B(_09774_),
    .C(_09882_),
    .X(_09883_));
 sky130_fd_sc_hd__a21o_1 _17345_ (.A1(_09773_),
    .A2(_09774_),
    .B1(_09882_),
    .X(_09884_));
 sky130_fd_sc_hd__or2b_2 _17346_ (.A(_09883_),
    .B_N(_09884_),
    .X(_09885_));
 sky130_fd_sc_hd__a21bo_1 _17347_ (.A1(_09759_),
    .A2(_09763_),
    .B1_N(_09757_),
    .X(_09886_));
 sky130_fd_sc_hd__xnor2_4 _17348_ (.A(_09885_),
    .B(_09886_),
    .Y(_09887_));
 sky130_fd_sc_hd__and2_1 _17349_ (.A(_09345_),
    .B(_09887_),
    .X(_09888_));
 sky130_fd_sc_hd__nand2_1 _17350_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .Y(_09889_));
 sky130_fd_sc_hd__or2_1 _17351_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .X(_09890_));
 sky130_fd_sc_hd__nand2_1 _17352_ (.A(_09766_),
    .B(_09770_),
    .Y(_09891_));
 sky130_fd_sc_hd__a21o_1 _17353_ (.A1(_09889_),
    .A2(_09890_),
    .B1(_09891_),
    .X(_09892_));
 sky130_fd_sc_hd__nand3_1 _17354_ (.A(_09889_),
    .B(_09890_),
    .C(_09891_),
    .Y(_09893_));
 sky130_fd_sc_hd__a31o_1 _17355_ (.A1(_09303_),
    .A2(_09892_),
    .A3(_09893_),
    .B1(_09282_),
    .X(_09894_));
 sky130_fd_sc_hd__o22a_1 _17356_ (.A1(\rbzero.wall_tracer.trackDistX[3] ),
    .A2(_09301_),
    .B1(_09888_),
    .B2(_09894_),
    .X(_00556_));
 sky130_fd_sc_hd__nor2_1 _17357_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .Y(_09895_));
 sky130_fd_sc_hd__and2_1 _17358_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .X(_09896_));
 sky130_fd_sc_hd__a21boi_1 _17359_ (.A1(_09890_),
    .A2(_09891_),
    .B1_N(_09889_),
    .Y(_09897_));
 sky130_fd_sc_hd__nor3_1 _17360_ (.A(_09895_),
    .B(_09896_),
    .C(_09897_),
    .Y(_09898_));
 sky130_fd_sc_hd__o21a_1 _17361_ (.A1(_09895_),
    .A2(_09896_),
    .B1(_09897_),
    .X(_09899_));
 sky130_fd_sc_hd__a31o_1 _17362_ (.A1(_09653_),
    .A2(_09655_),
    .A3(_09787_),
    .B1(_09785_),
    .X(_09900_));
 sky130_fd_sc_hd__nand2_1 _17363_ (.A(_09791_),
    .B(_09823_),
    .Y(_09901_));
 sky130_fd_sc_hd__or2b_1 _17364_ (.A(_09824_),
    .B_N(_09789_),
    .X(_09902_));
 sky130_fd_sc_hd__a21o_1 _17365_ (.A1(_09796_),
    .A2(_09806_),
    .B1(_09804_),
    .X(_09903_));
 sky130_fd_sc_hd__o31a_1 _17366_ (.A1(_07882_),
    .A2(_09115_),
    .A3(_09792_),
    .B1(_09793_),
    .X(_09904_));
 sky130_fd_sc_hd__inv_2 _17367_ (.A(_09904_),
    .Y(_09905_));
 sky130_fd_sc_hd__nand2_1 _17368_ (.A(_09903_),
    .B(_09905_),
    .Y(_09906_));
 sky130_fd_sc_hd__or2_1 _17369_ (.A(_09903_),
    .B(_09905_),
    .X(_09907_));
 sky130_fd_sc_hd__nand2_1 _17370_ (.A(_09906_),
    .B(_09907_),
    .Y(_09908_));
 sky130_fd_sc_hd__a21oi_1 _17371_ (.A1(_09901_),
    .A2(_09902_),
    .B1(_09908_),
    .Y(_09909_));
 sky130_fd_sc_hd__and3_1 _17372_ (.A(_09901_),
    .B(_09902_),
    .C(_09908_),
    .X(_09910_));
 sky130_fd_sc_hd__nor2_1 _17373_ (.A(_09909_),
    .B(_09910_),
    .Y(_09911_));
 sky130_fd_sc_hd__xnor2_2 _17374_ (.A(_09782_),
    .B(_09911_),
    .Y(_09912_));
 sky130_fd_sc_hd__a21o_1 _17375_ (.A1(_09807_),
    .A2(_09822_),
    .B1(_09820_),
    .X(_09913_));
 sky130_fd_sc_hd__or2_1 _17376_ (.A(_09828_),
    .B(_09844_),
    .X(_09914_));
 sky130_fd_sc_hd__o22a_1 _17377_ (.A1(_08890_),
    .A2(_08850_),
    .B1(_08979_),
    .B2(_08596_),
    .X(_09915_));
 sky130_fd_sc_hd__or4_1 _17378_ (.A(_08890_),
    .B(_08596_),
    .C(_08850_),
    .D(_08978_),
    .X(_09916_));
 sky130_fd_sc_hd__or2b_1 _17379_ (.A(_09915_),
    .B_N(_09916_),
    .X(_09917_));
 sky130_fd_sc_hd__nor2_1 _17380_ (.A(_08507_),
    .B(_09114_),
    .Y(_09918_));
 sky130_fd_sc_hd__xnor2_1 _17381_ (.A(_09917_),
    .B(_09918_),
    .Y(_09919_));
 sky130_fd_sc_hd__and3_1 _17382_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_03796_),
    .C(_08123_),
    .X(_09920_));
 sky130_fd_sc_hd__and3_1 _17383_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_03796_),
    .C(_08123_),
    .X(_09921_));
 sky130_fd_sc_hd__a21oi_1 _17384_ (.A1(_09018_),
    .A2(_08855_),
    .B1(_09921_),
    .Y(_09922_));
 sky130_fd_sc_hd__a21oi_1 _17385_ (.A1(_09797_),
    .A2(_09920_),
    .B1(_09922_),
    .Y(_09923_));
 sky130_fd_sc_hd__nor2_1 _17386_ (.A(_09022_),
    .B(_08723_),
    .Y(_09924_));
 sky130_fd_sc_hd__xnor2_1 _17387_ (.A(_09923_),
    .B(_09924_),
    .Y(_09925_));
 sky130_fd_sc_hd__o31a_1 _17388_ (.A1(_08890_),
    .A2(_08723_),
    .A3(_09798_),
    .B1(_09799_),
    .X(_09926_));
 sky130_fd_sc_hd__or2_1 _17389_ (.A(_09925_),
    .B(_09926_),
    .X(_09927_));
 sky130_fd_sc_hd__nand2_1 _17390_ (.A(_09925_),
    .B(_09926_),
    .Y(_09928_));
 sky130_fd_sc_hd__and2_1 _17391_ (.A(_09927_),
    .B(_09928_),
    .X(_09929_));
 sky130_fd_sc_hd__nand2_1 _17392_ (.A(_09919_),
    .B(_09929_),
    .Y(_09930_));
 sky130_fd_sc_hd__or2_1 _17393_ (.A(_09919_),
    .B(_09929_),
    .X(_09931_));
 sky130_fd_sc_hd__and2_1 _17394_ (.A(_09930_),
    .B(_09931_),
    .X(_09932_));
 sky130_fd_sc_hd__a21bo_1 _17395_ (.A1(_09811_),
    .A2(_09813_),
    .B1_N(_09810_),
    .X(_09933_));
 sky130_fd_sc_hd__a21bo_1 _17396_ (.A1(_09831_),
    .A2(_09834_),
    .B1_N(_09830_),
    .X(_09934_));
 sky130_fd_sc_hd__o22ai_1 _17397_ (.A1(_09833_),
    .A2(_07619_),
    .B1(_09571_),
    .B2(_08671_),
    .Y(_09935_));
 sky130_fd_sc_hd__or4_1 _17398_ (.A(_07472_),
    .B(_07618_),
    .C(_08732_),
    .D(_09571_),
    .X(_09936_));
 sky130_fd_sc_hd__nand2_1 _17399_ (.A(_09935_),
    .B(_09936_),
    .Y(_09937_));
 sky130_fd_sc_hd__nor2_1 _17400_ (.A(_09429_),
    .B(_07914_),
    .Y(_09938_));
 sky130_fd_sc_hd__xor2_1 _17401_ (.A(_09937_),
    .B(_09938_),
    .X(_09939_));
 sky130_fd_sc_hd__xnor2_1 _17402_ (.A(_09934_),
    .B(_09939_),
    .Y(_09940_));
 sky130_fd_sc_hd__xnor2_1 _17403_ (.A(_09933_),
    .B(_09940_),
    .Y(_09941_));
 sky130_fd_sc_hd__a21oi_1 _17404_ (.A1(_09808_),
    .A2(_09817_),
    .B1(_09815_),
    .Y(_09942_));
 sky130_fd_sc_hd__xor2_1 _17405_ (.A(_09941_),
    .B(_09942_),
    .X(_09943_));
 sky130_fd_sc_hd__nand2_1 _17406_ (.A(_09932_),
    .B(_09943_),
    .Y(_09944_));
 sky130_fd_sc_hd__or2_1 _17407_ (.A(_09932_),
    .B(_09943_),
    .X(_09945_));
 sky130_fd_sc_hd__nand2_1 _17408_ (.A(_09944_),
    .B(_09945_),
    .Y(_09946_));
 sky130_fd_sc_hd__a21o_1 _17409_ (.A1(_09914_),
    .A2(_09846_),
    .B1(_09946_),
    .X(_09947_));
 sky130_fd_sc_hd__nand3_1 _17410_ (.A(_09914_),
    .B(_09846_),
    .C(_09946_),
    .Y(_09948_));
 sky130_fd_sc_hd__nand2_1 _17411_ (.A(_09947_),
    .B(_09948_),
    .Y(_09949_));
 sky130_fd_sc_hd__xnor2_1 _17412_ (.A(_09913_),
    .B(_09949_),
    .Y(_09950_));
 sky130_fd_sc_hd__nor2_1 _17413_ (.A(_09840_),
    .B(_09842_),
    .Y(_09951_));
 sky130_fd_sc_hd__a21o_1 _17414_ (.A1(_09835_),
    .A2(_09843_),
    .B1(_09951_),
    .X(_09952_));
 sky130_fd_sc_hd__nor2_1 _17415_ (.A(_09850_),
    .B(_09854_),
    .Y(_09953_));
 sky130_fd_sc_hd__a21oi_1 _17416_ (.A1(_09849_),
    .A2(_09855_),
    .B1(_09953_),
    .Y(_09954_));
 sky130_fd_sc_hd__clkbuf_4 _17417_ (.A(_07663_),
    .X(_09955_));
 sky130_fd_sc_hd__or4_1 _17418_ (.A(_08594_),
    .B(_09428_),
    .C(_09955_),
    .D(_08780_),
    .X(_09956_));
 sky130_fd_sc_hd__a2bb2o_1 _17419_ (.A1_N(_09428_),
    .A2_N(_09955_),
    .B1(_08788_),
    .B2(_09163_),
    .X(_09957_));
 sky130_fd_sc_hd__nand2_1 _17420_ (.A(_09956_),
    .B(_09957_),
    .Y(_09958_));
 sky130_fd_sc_hd__nor2_1 _17421_ (.A(_07886_),
    .B(_09829_),
    .Y(_09959_));
 sky130_fd_sc_hd__xnor2_1 _17422_ (.A(_09958_),
    .B(_09959_),
    .Y(_09960_));
 sky130_fd_sc_hd__and2_1 _17423_ (.A(_07553_),
    .B(_09055_),
    .X(_09961_));
 sky130_fd_sc_hd__or2b_1 _17424_ (.A(_08240_),
    .B_N(_09055_),
    .X(_09962_));
 sky130_fd_sc_hd__nand2_1 _17425_ (.A(_08478_),
    .B(_08928_),
    .Y(_09963_));
 sky130_fd_sc_hd__nand2_1 _17426_ (.A(_07553_),
    .B(_09963_),
    .Y(_09964_));
 sky130_fd_sc_hd__a22o_1 _17427_ (.A1(_09836_),
    .A2(_09961_),
    .B1(_09962_),
    .B2(_09964_),
    .X(_09965_));
 sky130_fd_sc_hd__nor2_1 _17428_ (.A(_08760_),
    .B(_08917_),
    .Y(_09966_));
 sky130_fd_sc_hd__xor2_1 _17429_ (.A(_09965_),
    .B(_09966_),
    .X(_09967_));
 sky130_fd_sc_hd__buf_2 _17430_ (.A(_08760_),
    .X(_09968_));
 sky130_fd_sc_hd__o31a_1 _17431_ (.A1(_09968_),
    .A2(_08780_),
    .A3(_09838_),
    .B1(_09837_),
    .X(_09969_));
 sky130_fd_sc_hd__xor2_1 _17432_ (.A(_09967_),
    .B(_09969_),
    .X(_09970_));
 sky130_fd_sc_hd__xnor2_1 _17433_ (.A(_09960_),
    .B(_09970_),
    .Y(_09971_));
 sky130_fd_sc_hd__xor2_1 _17434_ (.A(_09954_),
    .B(_09971_),
    .X(_09972_));
 sky130_fd_sc_hd__xor2_1 _17435_ (.A(_09952_),
    .B(_09972_),
    .X(_09973_));
 sky130_fd_sc_hd__nor2_1 _17436_ (.A(_09449_),
    .B(_09603_),
    .Y(_09974_));
 sky130_fd_sc_hd__a22o_1 _17437_ (.A1(_09721_),
    .A2(_09974_),
    .B1(_09852_),
    .B2(_09853_),
    .X(_09975_));
 sky130_fd_sc_hd__o21a_4 _17438_ (.A1(_04939_),
    .A2(_09200_),
    .B1(_09731_),
    .X(_09976_));
 sky130_fd_sc_hd__o31ai_1 _17439_ (.A1(_09467_),
    .A2(_09728_),
    .A3(_09976_),
    .B1(_09465_),
    .Y(_09977_));
 sky130_fd_sc_hd__o21a_2 _17440_ (.A1(_04939_),
    .A2(_09051_),
    .B1(_09610_),
    .X(_09978_));
 sky130_fd_sc_hd__or3_1 _17441_ (.A(_09449_),
    .B(_09978_),
    .C(_09851_),
    .X(_09979_));
 sky130_fd_sc_hd__a22o_1 _17442_ (.A1(_08771_),
    .A2(_09607_),
    .B1(_09611_),
    .B2(_08046_),
    .X(_09980_));
 sky130_fd_sc_hd__or4bb_1 _17443_ (.A(_07858_),
    .B(_09463_),
    .C_N(_09979_),
    .D_N(_09980_),
    .X(_09981_));
 sky130_fd_sc_hd__a2bb2o_1 _17444_ (.A1_N(_09182_),
    .A2_N(_09463_),
    .B1(_09979_),
    .B2(_09980_),
    .X(_09982_));
 sky130_fd_sc_hd__nand3_1 _17445_ (.A(_09977_),
    .B(_09981_),
    .C(_09982_),
    .Y(_09983_));
 sky130_fd_sc_hd__a21o_1 _17446_ (.A1(_09981_),
    .A2(_09982_),
    .B1(_09977_),
    .X(_09984_));
 sky130_fd_sc_hd__and3_1 _17447_ (.A(_09975_),
    .B(_09983_),
    .C(_09984_),
    .X(_09985_));
 sky130_fd_sc_hd__a21oi_1 _17448_ (.A1(_09983_),
    .A2(_09984_),
    .B1(_09975_),
    .Y(_09986_));
 sky130_fd_sc_hd__nor2_1 _17449_ (.A(_07814_),
    .B(_09976_),
    .Y(_09987_));
 sky130_fd_sc_hd__mux2_1 _17450_ (.A0(_09987_),
    .A1(_07814_),
    .S(_09857_),
    .X(_09988_));
 sky130_fd_sc_hd__a21o_1 _17451_ (.A1(_09733_),
    .A2(_09735_),
    .B1(_09988_),
    .X(_09989_));
 sky130_fd_sc_hd__nand3_1 _17452_ (.A(_09733_),
    .B(_09735_),
    .C(_09988_),
    .Y(_09990_));
 sky130_fd_sc_hd__a21o_1 _17453_ (.A1(_09735_),
    .A2(_09858_),
    .B1(_09861_),
    .X(_09991_));
 sky130_fd_sc_hd__and3_1 _17454_ (.A(_09989_),
    .B(_09990_),
    .C(_09991_),
    .X(_09992_));
 sky130_fd_sc_hd__a21oi_1 _17455_ (.A1(_09989_),
    .A2(_09990_),
    .B1(_09991_),
    .Y(_09993_));
 sky130_fd_sc_hd__or4_1 _17456_ (.A(_09985_),
    .B(_09986_),
    .C(_09992_),
    .D(_09993_),
    .X(_09994_));
 sky130_fd_sc_hd__o22ai_1 _17457_ (.A1(_09985_),
    .A2(_09986_),
    .B1(_09992_),
    .B2(_09993_),
    .Y(_09995_));
 sky130_fd_sc_hd__a21o_1 _17458_ (.A1(_09856_),
    .A2(_09864_),
    .B1(_09863_),
    .X(_09996_));
 sky130_fd_sc_hd__nand3_1 _17459_ (.A(_09994_),
    .B(_09995_),
    .C(_09996_),
    .Y(_09997_));
 sky130_fd_sc_hd__a21o_1 _17460_ (.A1(_09994_),
    .A2(_09995_),
    .B1(_09996_),
    .X(_09998_));
 sky130_fd_sc_hd__and3_1 _17461_ (.A(_09973_),
    .B(_09997_),
    .C(_09998_),
    .X(_09999_));
 sky130_fd_sc_hd__a21oi_1 _17462_ (.A1(_09997_),
    .A2(_09998_),
    .B1(_09973_),
    .Y(_10000_));
 sky130_fd_sc_hd__or2_1 _17463_ (.A(_09999_),
    .B(_10000_),
    .X(_10001_));
 sky130_fd_sc_hd__and2_1 _17464_ (.A(_09866_),
    .B(_09868_),
    .X(_10002_));
 sky130_fd_sc_hd__a21oi_1 _17465_ (.A1(_09848_),
    .A2(_09869_),
    .B1(_10002_),
    .Y(_10003_));
 sky130_fd_sc_hd__xor2_1 _17466_ (.A(_10001_),
    .B(_10003_),
    .X(_10004_));
 sky130_fd_sc_hd__xnor2_1 _17467_ (.A(_09950_),
    .B(_10004_),
    .Y(_10005_));
 sky130_fd_sc_hd__nor2_1 _17468_ (.A(_09870_),
    .B(_09872_),
    .Y(_10006_));
 sky130_fd_sc_hd__a21oi_1 _17469_ (.A1(_09825_),
    .A2(_09873_),
    .B1(_10006_),
    .Y(_10007_));
 sky130_fd_sc_hd__nor2_1 _17470_ (.A(_10005_),
    .B(_10007_),
    .Y(_10008_));
 sky130_fd_sc_hd__and2_1 _17471_ (.A(_10005_),
    .B(_10007_),
    .X(_10009_));
 sky130_fd_sc_hd__nor2_1 _17472_ (.A(_10008_),
    .B(_10009_),
    .Y(_10010_));
 sky130_fd_sc_hd__xnor2_2 _17473_ (.A(_09912_),
    .B(_10010_),
    .Y(_10011_));
 sky130_fd_sc_hd__nor2_1 _17474_ (.A(_09874_),
    .B(_09876_),
    .Y(_10012_));
 sky130_fd_sc_hd__a21oi_1 _17475_ (.A1(_09788_),
    .A2(_09877_),
    .B1(_10012_),
    .Y(_10013_));
 sky130_fd_sc_hd__xnor2_1 _17476_ (.A(_10011_),
    .B(_10013_),
    .Y(_10014_));
 sky130_fd_sc_hd__xor2_1 _17477_ (.A(_09900_),
    .B(_10014_),
    .X(_10015_));
 sky130_fd_sc_hd__or2b_1 _17478_ (.A(_09881_),
    .B_N(_09776_),
    .X(_10016_));
 sky130_fd_sc_hd__o21a_1 _17479_ (.A1(_09878_),
    .A2(_09880_),
    .B1(_10016_),
    .X(_10017_));
 sky130_fd_sc_hd__nor2_1 _17480_ (.A(_10015_),
    .B(_10017_),
    .Y(_10018_));
 sky130_fd_sc_hd__and2_1 _17481_ (.A(_10015_),
    .B(_10017_),
    .X(_10019_));
 sky130_fd_sc_hd__or2_1 _17482_ (.A(_10018_),
    .B(_10019_),
    .X(_10020_));
 sky130_fd_sc_hd__a21o_1 _17483_ (.A1(_09757_),
    .A2(_09884_),
    .B1(_09883_),
    .X(_10021_));
 sky130_fd_sc_hd__nand2_1 _17484_ (.A(_09762_),
    .B(_10021_),
    .Y(_10022_));
 sky130_fd_sc_hd__a21o_1 _17485_ (.A1(_09369_),
    .A2(_09761_),
    .B1(_10022_),
    .X(_10023_));
 sky130_fd_sc_hd__a21oi_1 _17486_ (.A1(_09758_),
    .A2(_09884_),
    .B1(_09883_),
    .Y(_10024_));
 sky130_fd_sc_hd__nand2_1 _17487_ (.A(_10023_),
    .B(_10024_),
    .Y(_10025_));
 sky130_fd_sc_hd__or2_1 _17488_ (.A(_10020_),
    .B(_10025_),
    .X(_10026_));
 sky130_fd_sc_hd__nand2_1 _17489_ (.A(_04940_),
    .B(_10026_),
    .Y(_10027_));
 sky130_fd_sc_hd__a21o_1 _17490_ (.A1(_10020_),
    .A2(_10025_),
    .B1(_10027_),
    .X(_10028_));
 sky130_fd_sc_hd__o311a_1 _17491_ (.A1(_09345_),
    .A2(_09898_),
    .A3(_09899_),
    .B1(_09274_),
    .C1(_10028_),
    .X(_10029_));
 sky130_fd_sc_hd__a21oi_1 _17492_ (.A1(_07291_),
    .A2(_09283_),
    .B1(_10029_),
    .Y(_00557_));
 sky130_fd_sc_hd__nor2_1 _17493_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .Y(_10030_));
 sky130_fd_sc_hd__and2_1 _17494_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .X(_10031_));
 sky130_fd_sc_hd__o21ba_1 _17495_ (.A1(_09895_),
    .A2(_09897_),
    .B1_N(_09896_),
    .X(_10032_));
 sky130_fd_sc_hd__nor3_1 _17496_ (.A(_10030_),
    .B(_10031_),
    .C(_10032_),
    .Y(_10033_));
 sky130_fd_sc_hd__o21a_1 _17497_ (.A1(_10030_),
    .A2(_10031_),
    .B1(_10032_),
    .X(_10034_));
 sky130_fd_sc_hd__inv_2 _17498_ (.A(_10018_),
    .Y(_10035_));
 sky130_fd_sc_hd__or2_1 _17499_ (.A(_10011_),
    .B(_10013_),
    .X(_10036_));
 sky130_fd_sc_hd__or2b_1 _17500_ (.A(_10014_),
    .B_N(_09900_),
    .X(_10037_));
 sky130_fd_sc_hd__a31o_1 _17501_ (.A1(_09779_),
    .A2(_09781_),
    .A3(_09911_),
    .B1(_09909_),
    .X(_10038_));
 sky130_fd_sc_hd__or2b_1 _17502_ (.A(_09949_),
    .B_N(_09913_),
    .X(_10039_));
 sky130_fd_sc_hd__o31a_1 _17503_ (.A1(_08507_),
    .A2(_09115_),
    .A3(_09915_),
    .B1(_09916_),
    .X(_10040_));
 sky130_fd_sc_hd__a21oi_1 _17504_ (.A1(_09927_),
    .A2(_09930_),
    .B1(_10040_),
    .Y(_10041_));
 sky130_fd_sc_hd__and3_1 _17505_ (.A(_09927_),
    .B(_09930_),
    .C(_10040_),
    .X(_10042_));
 sky130_fd_sc_hd__or2_1 _17506_ (.A(_10041_),
    .B(_10042_),
    .X(_10043_));
 sky130_fd_sc_hd__a21oi_1 _17507_ (.A1(_09947_),
    .A2(_10039_),
    .B1(_10043_),
    .Y(_10044_));
 sky130_fd_sc_hd__and3_1 _17508_ (.A(_09947_),
    .B(_10039_),
    .C(_10043_),
    .X(_10045_));
 sky130_fd_sc_hd__nor2_1 _17509_ (.A(_10044_),
    .B(_10045_),
    .Y(_10046_));
 sky130_fd_sc_hd__xnor2_1 _17510_ (.A(_09906_),
    .B(_10046_),
    .Y(_10047_));
 sky130_fd_sc_hd__o21ai_1 _17511_ (.A1(_09941_),
    .A2(_09942_),
    .B1(_09944_),
    .Y(_10048_));
 sky130_fd_sc_hd__or2_1 _17512_ (.A(_09954_),
    .B(_09971_),
    .X(_10049_));
 sky130_fd_sc_hd__nand2_1 _17513_ (.A(_09952_),
    .B(_09972_),
    .Y(_10050_));
 sky130_fd_sc_hd__o22ai_1 _17514_ (.A1(_09022_),
    .A2(_08851_),
    .B1(_09373_),
    .B2(_08890_),
    .Y(_10051_));
 sky130_fd_sc_hd__or4_1 _17515_ (.A(_09022_),
    .B(_08890_),
    .C(_08851_),
    .D(_08979_),
    .X(_10052_));
 sky130_fd_sc_hd__nand2_1 _17516_ (.A(_10051_),
    .B(_10052_),
    .Y(_10053_));
 sky130_fd_sc_hd__and3_2 _17517_ (.A(_07420_),
    .B(_07421_),
    .C(_09389_),
    .X(_10054_));
 sky130_fd_sc_hd__xnor2_1 _17518_ (.A(_10053_),
    .B(_10054_),
    .Y(_10055_));
 sky130_fd_sc_hd__and2_2 _17519_ (.A(_07704_),
    .B(_07707_),
    .X(_10056_));
 sky130_fd_sc_hd__o21ba_1 _17520_ (.A1(_10056_),
    .A2(_08717_),
    .B1_N(_09920_),
    .X(_10057_));
 sky130_fd_sc_hd__nor2_1 _17521_ (.A(_10056_),
    .B(_08985_),
    .Y(_10058_));
 sky130_fd_sc_hd__nand2_1 _17522_ (.A(_09921_),
    .B(_10058_),
    .Y(_10059_));
 sky130_fd_sc_hd__or2b_1 _17523_ (.A(_10057_),
    .B_N(_10059_),
    .X(_10060_));
 sky130_fd_sc_hd__nor2_1 _17524_ (.A(_09684_),
    .B(_08723_),
    .Y(_10061_));
 sky130_fd_sc_hd__xor2_1 _17525_ (.A(_10060_),
    .B(_10061_),
    .X(_10062_));
 sky130_fd_sc_hd__nand2_1 _17526_ (.A(_09797_),
    .B(_09920_),
    .Y(_10063_));
 sky130_fd_sc_hd__o31a_1 _17527_ (.A1(_09022_),
    .A2(_08724_),
    .A3(_09922_),
    .B1(_10063_),
    .X(_10064_));
 sky130_fd_sc_hd__or2_1 _17528_ (.A(_10062_),
    .B(_10064_),
    .X(_10065_));
 sky130_fd_sc_hd__nand2_1 _17529_ (.A(_10062_),
    .B(_10064_),
    .Y(_10066_));
 sky130_fd_sc_hd__and2_1 _17530_ (.A(_10065_),
    .B(_10066_),
    .X(_10067_));
 sky130_fd_sc_hd__nand2_1 _17531_ (.A(_10055_),
    .B(_10067_),
    .Y(_10068_));
 sky130_fd_sc_hd__or2_1 _17532_ (.A(_10055_),
    .B(_10067_),
    .X(_10069_));
 sky130_fd_sc_hd__and2_1 _17533_ (.A(_10068_),
    .B(_10069_),
    .X(_10070_));
 sky130_fd_sc_hd__a21bo_1 _17534_ (.A1(_09935_),
    .A2(_09938_),
    .B1_N(_09936_),
    .X(_10071_));
 sky130_fd_sc_hd__a21bo_1 _17535_ (.A1(_09957_),
    .A2(_09959_),
    .B1_N(_09956_),
    .X(_10072_));
 sky130_fd_sc_hd__nor2_1 _17536_ (.A(_07472_),
    .B(_07618_),
    .Y(_10073_));
 sky130_fd_sc_hd__nor2_1 _17537_ (.A(_08732_),
    .B(_09829_),
    .Y(_10074_));
 sky130_fd_sc_hd__xnor2_1 _17538_ (.A(_10073_),
    .B(_10074_),
    .Y(_10075_));
 sky130_fd_sc_hd__or3_1 _17539_ (.A(_09571_),
    .B(_08735_),
    .C(_10075_),
    .X(_10076_));
 sky130_fd_sc_hd__o21ai_1 _17540_ (.A1(_09571_),
    .A2(_08735_),
    .B1(_10075_),
    .Y(_10077_));
 sky130_fd_sc_hd__nand2_1 _17541_ (.A(_10076_),
    .B(_10077_),
    .Y(_10078_));
 sky130_fd_sc_hd__xnor2_1 _17542_ (.A(_10072_),
    .B(_10078_),
    .Y(_10079_));
 sky130_fd_sc_hd__xnor2_1 _17543_ (.A(_10071_),
    .B(_10079_),
    .Y(_10080_));
 sky130_fd_sc_hd__and2b_1 _17544_ (.A_N(_09939_),
    .B(_09934_),
    .X(_10081_));
 sky130_fd_sc_hd__a21oi_1 _17545_ (.A1(_09933_),
    .A2(_09940_),
    .B1(_10081_),
    .Y(_10082_));
 sky130_fd_sc_hd__nor2_1 _17546_ (.A(_10080_),
    .B(_10082_),
    .Y(_10083_));
 sky130_fd_sc_hd__and2_1 _17547_ (.A(_10080_),
    .B(_10082_),
    .X(_10084_));
 sky130_fd_sc_hd__nor2_1 _17548_ (.A(_10083_),
    .B(_10084_),
    .Y(_10085_));
 sky130_fd_sc_hd__xnor2_1 _17549_ (.A(_10070_),
    .B(_10085_),
    .Y(_10086_));
 sky130_fd_sc_hd__a21o_1 _17550_ (.A1(_10049_),
    .A2(_10050_),
    .B1(_10086_),
    .X(_10087_));
 sky130_fd_sc_hd__nand3_1 _17551_ (.A(_10049_),
    .B(_10050_),
    .C(_10086_),
    .Y(_10088_));
 sky130_fd_sc_hd__nand2_1 _17552_ (.A(_10087_),
    .B(_10088_),
    .Y(_10089_));
 sky130_fd_sc_hd__xnor2_1 _17553_ (.A(_10048_),
    .B(_10089_),
    .Y(_10090_));
 sky130_fd_sc_hd__nor2_1 _17554_ (.A(_09967_),
    .B(_09969_),
    .Y(_10091_));
 sky130_fd_sc_hd__a21o_1 _17555_ (.A1(_09960_),
    .A2(_09970_),
    .B1(_10091_),
    .X(_10092_));
 sky130_fd_sc_hd__a21bo_1 _17556_ (.A1(_09975_),
    .A2(_09984_),
    .B1_N(_09983_),
    .X(_10093_));
 sky130_fd_sc_hd__or4_1 _17557_ (.A(_08594_),
    .B(_08595_),
    .C(_07840_),
    .D(_08917_),
    .X(_10094_));
 sky130_fd_sc_hd__clkbuf_4 _17558_ (.A(_07840_),
    .X(_10095_));
 sky130_fd_sc_hd__o22ai_1 _17559_ (.A1(_08595_),
    .A2(_10095_),
    .B1(_08917_),
    .B2(_08594_),
    .Y(_10096_));
 sky130_fd_sc_hd__nand2_1 _17560_ (.A(_10094_),
    .B(_10096_),
    .Y(_10097_));
 sky130_fd_sc_hd__nor2_1 _17561_ (.A(_07631_),
    .B(_09955_),
    .Y(_10098_));
 sky130_fd_sc_hd__xnor2_1 _17562_ (.A(_10097_),
    .B(_10098_),
    .Y(_10099_));
 sky130_fd_sc_hd__a21oi_1 _17563_ (.A1(_08787_),
    .A2(_09207_),
    .B1(_08240_),
    .Y(_10100_));
 sky130_fd_sc_hd__o32a_1 _17564_ (.A1(_08241_),
    .A2(_09463_),
    .A3(_09962_),
    .B1(_10100_),
    .B2(_09961_),
    .X(_10101_));
 sky130_fd_sc_hd__nor2_1 _17565_ (.A(_08760_),
    .B(_09451_),
    .Y(_10102_));
 sky130_fd_sc_hd__xnor2_1 _17566_ (.A(_10101_),
    .B(_10102_),
    .Y(_10103_));
 sky130_fd_sc_hd__nand2_1 _17567_ (.A(_09836_),
    .B(_09961_),
    .Y(_10104_));
 sky130_fd_sc_hd__o31a_1 _17568_ (.A1(_09968_),
    .A2(_08917_),
    .A3(_09965_),
    .B1(_10104_),
    .X(_10105_));
 sky130_fd_sc_hd__xor2_1 _17569_ (.A(_10103_),
    .B(_10105_),
    .X(_10106_));
 sky130_fd_sc_hd__xnor2_1 _17570_ (.A(_10099_),
    .B(_10106_),
    .Y(_10107_));
 sky130_fd_sc_hd__xor2_1 _17571_ (.A(_10093_),
    .B(_10107_),
    .X(_10108_));
 sky130_fd_sc_hd__xnor2_1 _17572_ (.A(_10092_),
    .B(_10108_),
    .Y(_10109_));
 sky130_fd_sc_hd__nand2_1 _17573_ (.A(_09979_),
    .B(_09981_),
    .Y(_10110_));
 sky130_fd_sc_hd__a21bo_4 _17574_ (.A1(_08779_),
    .A2(_09857_),
    .B1_N(_09465_),
    .X(_10111_));
 sky130_fd_sc_hd__a22o_1 _17575_ (.A1(_08771_),
    .A2(_09611_),
    .B1(_09732_),
    .B2(_08046_),
    .X(_10112_));
 sky130_fd_sc_hd__or4_1 _17576_ (.A(_08272_),
    .B(_09449_),
    .C(_09978_),
    .D(_09976_),
    .X(_10113_));
 sky130_fd_sc_hd__or4bb_1 _17577_ (.A(_07858_),
    .B(_09603_),
    .C_N(_10112_),
    .D_N(_10113_),
    .X(_10114_));
 sky130_fd_sc_hd__a2bb2o_1 _17578_ (.A1_N(_09182_),
    .A2_N(_09603_),
    .B1(_10112_),
    .B2(_10113_),
    .X(_10115_));
 sky130_fd_sc_hd__nand3_1 _17579_ (.A(_10111_),
    .B(_10114_),
    .C(_10115_),
    .Y(_10116_));
 sky130_fd_sc_hd__a21o_1 _17580_ (.A1(_10114_),
    .A2(_10115_),
    .B1(_10111_),
    .X(_10117_));
 sky130_fd_sc_hd__nand3_1 _17581_ (.A(_10110_),
    .B(_10116_),
    .C(_10117_),
    .Y(_10118_));
 sky130_fd_sc_hd__a21o_1 _17582_ (.A1(_10116_),
    .A2(_10117_),
    .B1(_10110_),
    .X(_10119_));
 sky130_fd_sc_hd__nand2_1 _17583_ (.A(_09861_),
    .B(_09988_),
    .Y(_10120_));
 sky130_fd_sc_hd__o21a_2 _17584_ (.A1(_09861_),
    .A2(_09989_),
    .B1(_10120_),
    .X(_10121_));
 sky130_fd_sc_hd__nand3_1 _17585_ (.A(_10118_),
    .B(_10119_),
    .C(_10121_),
    .Y(_10122_));
 sky130_fd_sc_hd__a21o_1 _17586_ (.A1(_10118_),
    .A2(_10119_),
    .B1(_10121_),
    .X(_10123_));
 sky130_fd_sc_hd__nand3_1 _17587_ (.A(_09989_),
    .B(_09990_),
    .C(_09991_),
    .Y(_10124_));
 sky130_fd_sc_hd__o31ai_1 _17588_ (.A1(_09985_),
    .A2(_09986_),
    .A3(_09993_),
    .B1(_10124_),
    .Y(_10125_));
 sky130_fd_sc_hd__nand3_1 _17589_ (.A(_10122_),
    .B(_10123_),
    .C(_10125_),
    .Y(_10126_));
 sky130_fd_sc_hd__a21o_1 _17590_ (.A1(_10122_),
    .A2(_10123_),
    .B1(_10125_),
    .X(_10127_));
 sky130_fd_sc_hd__and3_1 _17591_ (.A(_10109_),
    .B(_10126_),
    .C(_10127_),
    .X(_10128_));
 sky130_fd_sc_hd__a21oi_1 _17592_ (.A1(_10126_),
    .A2(_10127_),
    .B1(_10109_),
    .Y(_10129_));
 sky130_fd_sc_hd__or2_1 _17593_ (.A(_10128_),
    .B(_10129_),
    .X(_10130_));
 sky130_fd_sc_hd__a21boi_1 _17594_ (.A1(_09973_),
    .A2(_09998_),
    .B1_N(_09997_),
    .Y(_10131_));
 sky130_fd_sc_hd__xor2_1 _17595_ (.A(_10130_),
    .B(_10131_),
    .X(_10132_));
 sky130_fd_sc_hd__xnor2_1 _17596_ (.A(_10090_),
    .B(_10132_),
    .Y(_10133_));
 sky130_fd_sc_hd__nor2_1 _17597_ (.A(_10001_),
    .B(_10003_),
    .Y(_10134_));
 sky130_fd_sc_hd__a21oi_1 _17598_ (.A1(_09950_),
    .A2(_10004_),
    .B1(_10134_),
    .Y(_10135_));
 sky130_fd_sc_hd__nor2_1 _17599_ (.A(_10133_),
    .B(_10135_),
    .Y(_10136_));
 sky130_fd_sc_hd__and2_1 _17600_ (.A(_10133_),
    .B(_10135_),
    .X(_10137_));
 sky130_fd_sc_hd__nor2_1 _17601_ (.A(_10136_),
    .B(_10137_),
    .Y(_10138_));
 sky130_fd_sc_hd__xnor2_1 _17602_ (.A(_10047_),
    .B(_10138_),
    .Y(_10139_));
 sky130_fd_sc_hd__a21oi_1 _17603_ (.A1(_09912_),
    .A2(_10010_),
    .B1(_10008_),
    .Y(_10140_));
 sky130_fd_sc_hd__xnor2_1 _17604_ (.A(_10139_),
    .B(_10140_),
    .Y(_10141_));
 sky130_fd_sc_hd__xor2_2 _17605_ (.A(_10038_),
    .B(_10141_),
    .X(_10142_));
 sky130_fd_sc_hd__a21oi_1 _17606_ (.A1(_10036_),
    .A2(_10037_),
    .B1(_10142_),
    .Y(_10143_));
 sky130_fd_sc_hd__nand3_1 _17607_ (.A(_10036_),
    .B(_10037_),
    .C(_10142_),
    .Y(_10144_));
 sky130_fd_sc_hd__or2b_1 _17608_ (.A(_10143_),
    .B_N(_10144_),
    .X(_10145_));
 sky130_fd_sc_hd__and3_1 _17609_ (.A(_10035_),
    .B(_10026_),
    .C(_10145_),
    .X(_10146_));
 sky130_fd_sc_hd__a21o_1 _17610_ (.A1(_10035_),
    .A2(_10026_),
    .B1(_10145_),
    .X(_10147_));
 sky130_fd_sc_hd__or3b_2 _17611_ (.A(_03797_),
    .B(_10146_),
    .C_N(_10147_),
    .X(_10148_));
 sky130_fd_sc_hd__o311a_1 _17612_ (.A1(_09345_),
    .A2(_10033_),
    .A3(_10034_),
    .B1(_09274_),
    .C1(_10148_),
    .X(_10149_));
 sky130_fd_sc_hd__a21oi_1 _17613_ (.A1(_07294_),
    .A2(_09283_),
    .B1(_10149_),
    .Y(_00558_));
 sky130_fd_sc_hd__or2_1 _17614_ (.A(_10139_),
    .B(_10140_),
    .X(_10150_));
 sky130_fd_sc_hd__or2b_1 _17615_ (.A(_10141_),
    .B_N(_10038_),
    .X(_10151_));
 sky130_fd_sc_hd__a31o_1 _17616_ (.A1(_09903_),
    .A2(_09905_),
    .A3(_10046_),
    .B1(_10044_),
    .X(_10152_));
 sky130_fd_sc_hd__or2b_1 _17617_ (.A(_10089_),
    .B_N(_10048_),
    .X(_10153_));
 sky130_fd_sc_hd__a21boi_1 _17618_ (.A1(_10051_),
    .A2(_10054_),
    .B1_N(_10052_),
    .Y(_10154_));
 sky130_fd_sc_hd__a21o_1 _17619_ (.A1(_10065_),
    .A2(_10068_),
    .B1(_10154_),
    .X(_10155_));
 sky130_fd_sc_hd__nand3_1 _17620_ (.A(_10065_),
    .B(_10068_),
    .C(_10154_),
    .Y(_10156_));
 sky130_fd_sc_hd__nand2_1 _17621_ (.A(_10155_),
    .B(_10156_),
    .Y(_10157_));
 sky130_fd_sc_hd__a21oi_1 _17622_ (.A1(_10087_),
    .A2(_10153_),
    .B1(_10157_),
    .Y(_10158_));
 sky130_fd_sc_hd__and3_1 _17623_ (.A(_10087_),
    .B(_10153_),
    .C(_10157_),
    .X(_10159_));
 sky130_fd_sc_hd__nor2_1 _17624_ (.A(_10158_),
    .B(_10159_),
    .Y(_10160_));
 sky130_fd_sc_hd__xor2_1 _17625_ (.A(_10041_),
    .B(_10160_),
    .X(_10161_));
 sky130_fd_sc_hd__a21o_1 _17626_ (.A1(_10070_),
    .A2(_10085_),
    .B1(_10083_),
    .X(_10162_));
 sky130_fd_sc_hd__or2b_1 _17627_ (.A(_10107_),
    .B_N(_10093_),
    .X(_10163_));
 sky130_fd_sc_hd__or2b_1 _17628_ (.A(_10108_),
    .B_N(_10092_),
    .X(_10164_));
 sky130_fd_sc_hd__o22a_1 _17629_ (.A1(_09684_),
    .A2(_08851_),
    .B1(_08979_),
    .B2(_09022_),
    .X(_10165_));
 sky130_fd_sc_hd__or4_1 _17630_ (.A(_09684_),
    .B(_09022_),
    .C(_08850_),
    .D(_08978_),
    .X(_10166_));
 sky130_fd_sc_hd__or2b_1 _17631_ (.A(_10165_),
    .B_N(_10166_),
    .X(_10167_));
 sky130_fd_sc_hd__nor2_1 _17632_ (.A(_08750_),
    .B(_09114_),
    .Y(_10168_));
 sky130_fd_sc_hd__xnor2_1 _17633_ (.A(_10167_),
    .B(_10168_),
    .Y(_10169_));
 sky130_fd_sc_hd__nor2_1 _17634_ (.A(_09571_),
    .B(_08717_),
    .Y(_10170_));
 sky130_fd_sc_hd__xnor2_1 _17635_ (.A(_10058_),
    .B(_10170_),
    .Y(_10171_));
 sky130_fd_sc_hd__or2_1 _17636_ (.A(_09166_),
    .B(_08723_),
    .X(_10172_));
 sky130_fd_sc_hd__xnor2_1 _17637_ (.A(_10171_),
    .B(_10172_),
    .Y(_10173_));
 sky130_fd_sc_hd__o31a_1 _17638_ (.A1(_09684_),
    .A2(_08723_),
    .A3(_10057_),
    .B1(_10059_),
    .X(_10174_));
 sky130_fd_sc_hd__or2_1 _17639_ (.A(_10173_),
    .B(_10174_),
    .X(_01424_));
 sky130_fd_sc_hd__nand2_1 _17640_ (.A(_10173_),
    .B(_10174_),
    .Y(_01425_));
 sky130_fd_sc_hd__and2_1 _17641_ (.A(_01424_),
    .B(_01425_),
    .X(_01426_));
 sky130_fd_sc_hd__nand2_1 _17642_ (.A(_10169_),
    .B(_01426_),
    .Y(_01427_));
 sky130_fd_sc_hd__or2_1 _17643_ (.A(_10169_),
    .B(_01426_),
    .X(_01428_));
 sky130_fd_sc_hd__and2_1 _17644_ (.A(_01427_),
    .B(_01428_),
    .X(_01429_));
 sky130_fd_sc_hd__a21bo_1 _17645_ (.A1(_10073_),
    .A2(_10074_),
    .B1_N(_10076_),
    .X(_01430_));
 sky130_fd_sc_hd__a21bo_1 _17646_ (.A1(_10096_),
    .A2(_10098_),
    .B1_N(_10094_),
    .X(_01431_));
 sky130_fd_sc_hd__a2bb2o_1 _17647_ (.A1_N(_07619_),
    .A2_N(_07663_),
    .B1(_08536_),
    .B2(_07651_),
    .X(_01432_));
 sky130_fd_sc_hd__or3b_1 _17648_ (.A(_07618_),
    .B(_07663_),
    .C_N(_10074_),
    .X(_01433_));
 sky130_fd_sc_hd__nand2_1 _17649_ (.A(_01432_),
    .B(_01433_),
    .Y(_01434_));
 sky130_fd_sc_hd__nor2_1 _17650_ (.A(_09833_),
    .B(_07914_),
    .Y(_01435_));
 sky130_fd_sc_hd__xnor2_1 _17651_ (.A(_01434_),
    .B(_01435_),
    .Y(_01436_));
 sky130_fd_sc_hd__xor2_1 _17652_ (.A(_01431_),
    .B(_01436_),
    .X(_01437_));
 sky130_fd_sc_hd__xnor2_1 _17653_ (.A(_01430_),
    .B(_01437_),
    .Y(_01438_));
 sky130_fd_sc_hd__and2b_1 _17654_ (.A_N(_10078_),
    .B(_10072_),
    .X(_01439_));
 sky130_fd_sc_hd__a21oi_1 _17655_ (.A1(_10071_),
    .A2(_10079_),
    .B1(_01439_),
    .Y(_01440_));
 sky130_fd_sc_hd__nor2_1 _17656_ (.A(_01438_),
    .B(_01440_),
    .Y(_01441_));
 sky130_fd_sc_hd__and2_1 _17657_ (.A(_01438_),
    .B(_01440_),
    .X(_01442_));
 sky130_fd_sc_hd__nor2_1 _17658_ (.A(_01441_),
    .B(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hd__xnor2_1 _17659_ (.A(_01429_),
    .B(_01443_),
    .Y(_01444_));
 sky130_fd_sc_hd__a21o_1 _17660_ (.A1(_10163_),
    .A2(_10164_),
    .B1(_01444_),
    .X(_01445_));
 sky130_fd_sc_hd__nand3_1 _17661_ (.A(_10163_),
    .B(_10164_),
    .C(_01444_),
    .Y(_01446_));
 sky130_fd_sc_hd__nand2_1 _17662_ (.A(_01445_),
    .B(_01446_),
    .Y(_01447_));
 sky130_fd_sc_hd__xnor2_1 _17663_ (.A(_10162_),
    .B(_01447_),
    .Y(_01448_));
 sky130_fd_sc_hd__nor2_1 _17664_ (.A(_10103_),
    .B(_10105_),
    .Y(_01449_));
 sky130_fd_sc_hd__a21o_1 _17665_ (.A1(_10099_),
    .A2(_10106_),
    .B1(_01449_),
    .X(_01450_));
 sky130_fd_sc_hd__nand2_1 _17666_ (.A(_10116_),
    .B(_10118_),
    .Y(_01451_));
 sky130_fd_sc_hd__or4_1 _17667_ (.A(_08067_),
    .B(_09428_),
    .C(_07827_),
    .D(_09451_),
    .X(_01452_));
 sky130_fd_sc_hd__a2bb2o_1 _17668_ (.A1_N(_09428_),
    .A2_N(_07827_),
    .B1(_09963_),
    .B2(_09163_),
    .X(_01453_));
 sky130_fd_sc_hd__nand2_1 _17669_ (.A(_01452_),
    .B(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__or3_1 _17670_ (.A(_07886_),
    .B(_10095_),
    .C(_01454_),
    .X(_01455_));
 sky130_fd_sc_hd__o21ai_1 _17671_ (.A1(_07886_),
    .A2(_10095_),
    .B1(_01454_),
    .Y(_01456_));
 sky130_fd_sc_hd__and2_1 _17672_ (.A(_01455_),
    .B(_01456_),
    .X(_01457_));
 sky130_fd_sc_hd__a21o_1 _17673_ (.A1(_08923_),
    .A2(_09470_),
    .B1(_08240_),
    .X(_01458_));
 sky130_fd_sc_hd__o21a_1 _17674_ (.A1(_08241_),
    .A2(_09462_),
    .B1(_01458_),
    .X(_01459_));
 sky130_fd_sc_hd__a21oi_1 _17675_ (.A1(_08923_),
    .A2(_09470_),
    .B1(_08241_),
    .Y(_01460_));
 sky130_fd_sc_hd__nand2_1 _17676_ (.A(_10100_),
    .B(_01460_),
    .Y(_01461_));
 sky130_fd_sc_hd__and2b_1 _17677_ (.A_N(_01459_),
    .B(_01461_),
    .X(_01462_));
 sky130_fd_sc_hd__nor2_1 _17678_ (.A(_09968_),
    .B(_09197_),
    .Y(_01463_));
 sky130_fd_sc_hd__xnor2_1 _17679_ (.A(_01462_),
    .B(_01463_),
    .Y(_01464_));
 sky130_fd_sc_hd__nand2_1 _17680_ (.A(_10101_),
    .B(_10102_),
    .Y(_01465_));
 sky130_fd_sc_hd__o31a_1 _17681_ (.A1(_08241_),
    .A2(_09463_),
    .A3(_09962_),
    .B1(_01465_),
    .X(_01466_));
 sky130_fd_sc_hd__xor2_1 _17682_ (.A(_01464_),
    .B(_01466_),
    .X(_01467_));
 sky130_fd_sc_hd__xor2_1 _17683_ (.A(_01457_),
    .B(_01467_),
    .X(_01468_));
 sky130_fd_sc_hd__xnor2_1 _17684_ (.A(_01451_),
    .B(_01468_),
    .Y(_01469_));
 sky130_fd_sc_hd__xnor2_1 _17685_ (.A(_01450_),
    .B(_01469_),
    .Y(_01470_));
 sky130_fd_sc_hd__nand2_1 _17686_ (.A(_10113_),
    .B(_10114_),
    .Y(_01471_));
 sky130_fd_sc_hd__or3_2 _17687_ (.A(_08272_),
    .B(_09449_),
    .C(_09976_),
    .X(_01472_));
 sky130_fd_sc_hd__a21oi_1 _17688_ (.A1(_08272_),
    .A2(_09449_),
    .B1(_09976_),
    .Y(_01473_));
 sky130_fd_sc_hd__or4bb_1 _17689_ (.A(_09182_),
    .B(_09978_),
    .C_N(_01472_),
    .D_N(_01473_),
    .X(_01474_));
 sky130_fd_sc_hd__a2bb2o_1 _17690_ (.A1_N(_09182_),
    .A2_N(_09978_),
    .B1(_01472_),
    .B2(_01473_),
    .X(_01475_));
 sky130_fd_sc_hd__nand3_1 _17691_ (.A(_10111_),
    .B(_01474_),
    .C(_01475_),
    .Y(_01476_));
 sky130_fd_sc_hd__a21o_1 _17692_ (.A1(_01474_),
    .A2(_01475_),
    .B1(_10111_),
    .X(_01477_));
 sky130_fd_sc_hd__nand3_1 _17693_ (.A(_01471_),
    .B(_01476_),
    .C(_01477_),
    .Y(_01478_));
 sky130_fd_sc_hd__a21o_1 _17694_ (.A1(_01476_),
    .A2(_01477_),
    .B1(_01471_),
    .X(_01479_));
 sky130_fd_sc_hd__and3_1 _17695_ (.A(_10121_),
    .B(_01478_),
    .C(_01479_),
    .X(_01480_));
 sky130_fd_sc_hd__a21oi_1 _17696_ (.A1(_01478_),
    .A2(_01479_),
    .B1(_10121_),
    .Y(_01481_));
 sky130_fd_sc_hd__a211oi_1 _17697_ (.A1(_10120_),
    .A2(_10122_),
    .B1(_01480_),
    .C1(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__o211a_1 _17698_ (.A1(_01480_),
    .A2(_01481_),
    .B1(_10120_),
    .C1(_10122_),
    .X(_01483_));
 sky130_fd_sc_hd__nor2_1 _17699_ (.A(_01482_),
    .B(_01483_),
    .Y(_01484_));
 sky130_fd_sc_hd__xnor2_1 _17700_ (.A(_01470_),
    .B(_01484_),
    .Y(_01485_));
 sky130_fd_sc_hd__a21boi_1 _17701_ (.A1(_10109_),
    .A2(_10127_),
    .B1_N(_10126_),
    .Y(_01486_));
 sky130_fd_sc_hd__xor2_1 _17702_ (.A(_01485_),
    .B(_01486_),
    .X(_01487_));
 sky130_fd_sc_hd__xnor2_1 _17703_ (.A(_01448_),
    .B(_01487_),
    .Y(_01488_));
 sky130_fd_sc_hd__nor2_1 _17704_ (.A(_10130_),
    .B(_10131_),
    .Y(_01489_));
 sky130_fd_sc_hd__a21oi_1 _17705_ (.A1(_10090_),
    .A2(_10132_),
    .B1(_01489_),
    .Y(_01490_));
 sky130_fd_sc_hd__nor2_1 _17706_ (.A(_01488_),
    .B(_01490_),
    .Y(_01491_));
 sky130_fd_sc_hd__nand2_1 _17707_ (.A(_01488_),
    .B(_01490_),
    .Y(_01492_));
 sky130_fd_sc_hd__and2b_1 _17708_ (.A_N(_01491_),
    .B(_01492_),
    .X(_01493_));
 sky130_fd_sc_hd__xnor2_1 _17709_ (.A(_10161_),
    .B(_01493_),
    .Y(_01494_));
 sky130_fd_sc_hd__a21oi_1 _17710_ (.A1(_10047_),
    .A2(_10138_),
    .B1(_10136_),
    .Y(_01495_));
 sky130_fd_sc_hd__xnor2_1 _17711_ (.A(_01494_),
    .B(_01495_),
    .Y(_01496_));
 sky130_fd_sc_hd__xor2_1 _17712_ (.A(_10152_),
    .B(_01496_),
    .X(_01497_));
 sky130_fd_sc_hd__a21o_2 _17713_ (.A1(_10150_),
    .A2(_10151_),
    .B1(_01497_),
    .X(_01498_));
 sky130_fd_sc_hd__nand3_1 _17714_ (.A(_10150_),
    .B(_10151_),
    .C(_01497_),
    .Y(_01499_));
 sky130_fd_sc_hd__nand2_2 _17715_ (.A(_01498_),
    .B(_01499_),
    .Y(_01500_));
 sky130_fd_sc_hd__nor2_1 _17716_ (.A(_10020_),
    .B(_10145_),
    .Y(_01501_));
 sky130_fd_sc_hd__a21o_1 _17717_ (.A1(_10018_),
    .A2(_10144_),
    .B1(_10143_),
    .X(_01502_));
 sky130_fd_sc_hd__a31oi_1 _17718_ (.A1(_10023_),
    .A2(_10024_),
    .A3(_01501_),
    .B1(_01502_),
    .Y(_01503_));
 sky130_fd_sc_hd__or2_1 _17719_ (.A(_01500_),
    .B(_01503_),
    .X(_01504_));
 sky130_fd_sc_hd__nand2_1 _17720_ (.A(_09345_),
    .B(_01504_),
    .Y(_01505_));
 sky130_fd_sc_hd__a21oi_2 _17721_ (.A1(_01500_),
    .A2(_01503_),
    .B1(_01505_),
    .Y(_01506_));
 sky130_fd_sc_hd__nor2_1 _17722_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .Y(_01507_));
 sky130_fd_sc_hd__and2_1 _17723_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .X(_01508_));
 sky130_fd_sc_hd__o21ba_1 _17724_ (.A1(_10030_),
    .A2(_10032_),
    .B1_N(_10031_),
    .X(_01509_));
 sky130_fd_sc_hd__or3_1 _17725_ (.A(_01507_),
    .B(_01508_),
    .C(_01509_),
    .X(_01510_));
 sky130_fd_sc_hd__o21ai_1 _17726_ (.A1(_01507_),
    .A2(_01508_),
    .B1(_01509_),
    .Y(_01511_));
 sky130_fd_sc_hd__a31o_1 _17727_ (.A1(_09303_),
    .A2(_01510_),
    .A3(_01511_),
    .B1(_09282_),
    .X(_01512_));
 sky130_fd_sc_hd__o22a_1 _17728_ (.A1(\rbzero.wall_tracer.trackDistX[6] ),
    .A2(_09275_),
    .B1(_01506_),
    .B2(_01512_),
    .X(_00559_));
 sky130_fd_sc_hd__or2_1 _17729_ (.A(_01494_),
    .B(_01495_),
    .X(_01513_));
 sky130_fd_sc_hd__or2b_1 _17730_ (.A(_01496_),
    .B_N(_10152_),
    .X(_01514_));
 sky130_fd_sc_hd__a21o_1 _17731_ (.A1(_10041_),
    .A2(_10160_),
    .B1(_10158_),
    .X(_01515_));
 sky130_fd_sc_hd__or2b_1 _17732_ (.A(_01447_),
    .B_N(_10162_),
    .X(_01516_));
 sky130_fd_sc_hd__o31a_1 _17733_ (.A1(_08750_),
    .A2(_09115_),
    .A3(_10165_),
    .B1(_10166_),
    .X(_01517_));
 sky130_fd_sc_hd__a21o_1 _17734_ (.A1(_01424_),
    .A2(_01427_),
    .B1(_01517_),
    .X(_01518_));
 sky130_fd_sc_hd__nand3_1 _17735_ (.A(_01424_),
    .B(_01427_),
    .C(_01517_),
    .Y(_01519_));
 sky130_fd_sc_hd__nand2_1 _17736_ (.A(_01518_),
    .B(_01519_),
    .Y(_01520_));
 sky130_fd_sc_hd__a21o_1 _17737_ (.A1(_01445_),
    .A2(_01516_),
    .B1(_01520_),
    .X(_01521_));
 sky130_fd_sc_hd__nand3_1 _17738_ (.A(_01445_),
    .B(_01516_),
    .C(_01520_),
    .Y(_01522_));
 sky130_fd_sc_hd__and2_1 _17739_ (.A(_01521_),
    .B(_01522_),
    .X(_01523_));
 sky130_fd_sc_hd__xnor2_1 _17740_ (.A(_10155_),
    .B(_01523_),
    .Y(_01524_));
 sky130_fd_sc_hd__a21o_1 _17741_ (.A1(_01429_),
    .A2(_01443_),
    .B1(_01441_),
    .X(_01525_));
 sky130_fd_sc_hd__and2b_1 _17742_ (.A_N(_01469_),
    .B(_01450_),
    .X(_01526_));
 sky130_fd_sc_hd__a21o_1 _17743_ (.A1(_01451_),
    .A2(_01468_),
    .B1(_01526_),
    .X(_01527_));
 sky130_fd_sc_hd__nor2_1 _17744_ (.A(_09684_),
    .B(_08852_),
    .Y(_01528_));
 sky130_fd_sc_hd__nor2_1 _17745_ (.A(_09166_),
    .B(_08979_),
    .Y(_01529_));
 sky130_fd_sc_hd__o22a_1 _17746_ (.A1(_09166_),
    .A2(_08851_),
    .B1(_08979_),
    .B2(_09684_),
    .X(_01530_));
 sky130_fd_sc_hd__a21o_1 _17747_ (.A1(_01528_),
    .A2(_01529_),
    .B1(_01530_),
    .X(_01531_));
 sky130_fd_sc_hd__nor2_1 _17748_ (.A(_08135_),
    .B(_09115_),
    .Y(_01532_));
 sky130_fd_sc_hd__xnor2_1 _17749_ (.A(_01531_),
    .B(_01532_),
    .Y(_01533_));
 sky130_fd_sc_hd__o22a_1 _17750_ (.A1(_09833_),
    .A2(_08531_),
    .B1(_08985_),
    .B2(_09571_),
    .X(_01534_));
 sky130_fd_sc_hd__or2_1 _17751_ (.A(_07472_),
    .B(_08663_),
    .X(_01535_));
 sky130_fd_sc_hd__or3_1 _17752_ (.A(_09571_),
    .B(_08717_),
    .C(_01535_),
    .X(_01536_));
 sky130_fd_sc_hd__and2b_1 _17753_ (.A_N(_01534_),
    .B(_01536_),
    .X(_01537_));
 sky130_fd_sc_hd__nor2_1 _17754_ (.A(_10056_),
    .B(_08724_),
    .Y(_01538_));
 sky130_fd_sc_hd__xnor2_1 _17755_ (.A(_01537_),
    .B(_01538_),
    .Y(_01539_));
 sky130_fd_sc_hd__nand2_1 _17756_ (.A(_10058_),
    .B(_10170_),
    .Y(_01540_));
 sky130_fd_sc_hd__o31a_1 _17757_ (.A1(_09166_),
    .A2(_08724_),
    .A3(_10171_),
    .B1(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__or2_1 _17758_ (.A(_01539_),
    .B(_01541_),
    .X(_01542_));
 sky130_fd_sc_hd__nand2_1 _17759_ (.A(_01539_),
    .B(_01541_),
    .Y(_01543_));
 sky130_fd_sc_hd__and2_1 _17760_ (.A(_01542_),
    .B(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__nand2_1 _17761_ (.A(_01533_),
    .B(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hd__or2_1 _17762_ (.A(_01533_),
    .B(_01544_),
    .X(_01546_));
 sky130_fd_sc_hd__and2_1 _17763_ (.A(_01545_),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__a21bo_1 _17764_ (.A1(_01432_),
    .A2(_01435_),
    .B1_N(_01433_),
    .X(_01548_));
 sky130_fd_sc_hd__nand2_1 _17765_ (.A(_01452_),
    .B(_01455_),
    .Y(_01549_));
 sky130_fd_sc_hd__or4_1 _17766_ (.A(_07618_),
    .B(_08732_),
    .C(_09955_),
    .D(_10095_),
    .X(_01550_));
 sky130_fd_sc_hd__o22ai_1 _17767_ (.A1(_07618_),
    .A2(_09955_),
    .B1(_10095_),
    .B2(_08732_),
    .Y(_01551_));
 sky130_fd_sc_hd__nand2_1 _17768_ (.A(_01550_),
    .B(_01551_),
    .Y(_01552_));
 sky130_fd_sc_hd__nor2_1 _17769_ (.A(_09829_),
    .B(_08735_),
    .Y(_01553_));
 sky130_fd_sc_hd__xor2_1 _17770_ (.A(_01552_),
    .B(_01553_),
    .X(_01554_));
 sky130_fd_sc_hd__xnor2_1 _17771_ (.A(_01549_),
    .B(_01554_),
    .Y(_01555_));
 sky130_fd_sc_hd__xnor2_1 _17772_ (.A(_01548_),
    .B(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__and2_1 _17773_ (.A(_01431_),
    .B(_01436_),
    .X(_01557_));
 sky130_fd_sc_hd__a21oi_1 _17774_ (.A1(_01430_),
    .A2(_01437_),
    .B1(_01557_),
    .Y(_01558_));
 sky130_fd_sc_hd__nor2_1 _17775_ (.A(_01556_),
    .B(_01558_),
    .Y(_01559_));
 sky130_fd_sc_hd__nand2_1 _17776_ (.A(_01556_),
    .B(_01558_),
    .Y(_01560_));
 sky130_fd_sc_hd__and2b_1 _17777_ (.A_N(_01559_),
    .B(_01560_),
    .X(_01561_));
 sky130_fd_sc_hd__xnor2_1 _17778_ (.A(_01547_),
    .B(_01561_),
    .Y(_01562_));
 sky130_fd_sc_hd__xor2_1 _17779_ (.A(_01527_),
    .B(_01562_),
    .X(_01563_));
 sky130_fd_sc_hd__xnor2_2 _17780_ (.A(_01525_),
    .B(_01563_),
    .Y(_01564_));
 sky130_fd_sc_hd__nor2_1 _17781_ (.A(_01464_),
    .B(_01466_),
    .Y(_01565_));
 sky130_fd_sc_hd__a21o_1 _17782_ (.A1(_01457_),
    .A2(_01467_),
    .B1(_01565_),
    .X(_01566_));
 sky130_fd_sc_hd__nand2_1 _17783_ (.A(_01476_),
    .B(_01478_),
    .Y(_01567_));
 sky130_fd_sc_hd__or4_1 _17784_ (.A(_08067_),
    .B(_08595_),
    .C(_08645_),
    .D(_09197_),
    .X(_01568_));
 sky130_fd_sc_hd__a2bb2o_1 _17785_ (.A1_N(_08595_),
    .A2_N(_08645_),
    .B1(_09055_),
    .B2(_09163_),
    .X(_01569_));
 sky130_fd_sc_hd__nand2_1 _17786_ (.A(_01568_),
    .B(_01569_),
    .Y(_01570_));
 sky130_fd_sc_hd__or3_1 _17787_ (.A(_07631_),
    .B(_07827_),
    .C(_01570_),
    .X(_01571_));
 sky130_fd_sc_hd__o21ai_1 _17788_ (.A1(_07631_),
    .A2(_07827_),
    .B1(_01570_),
    .Y(_01572_));
 sky130_fd_sc_hd__and2_1 _17789_ (.A(_01571_),
    .B(_01572_),
    .X(_01573_));
 sky130_fd_sc_hd__nand2_1 _17790_ (.A(_07553_),
    .B(_09611_),
    .Y(_01574_));
 sky130_fd_sc_hd__o21bai_1 _17791_ (.A1(_08240_),
    .A2(_09978_),
    .B1_N(_01460_),
    .Y(_01575_));
 sky130_fd_sc_hd__o21ai_1 _17792_ (.A1(_01458_),
    .A2(_01574_),
    .B1(_01575_),
    .Y(_01576_));
 sky130_fd_sc_hd__nor2_1 _17793_ (.A(_09968_),
    .B(_09463_),
    .Y(_01577_));
 sky130_fd_sc_hd__xor2_1 _17794_ (.A(_01576_),
    .B(_01577_),
    .X(_01578_));
 sky130_fd_sc_hd__o31a_1 _17795_ (.A1(_09968_),
    .A2(_09197_),
    .A3(_01459_),
    .B1(_01461_),
    .X(_01579_));
 sky130_fd_sc_hd__xor2_1 _17796_ (.A(_01578_),
    .B(_01579_),
    .X(_01580_));
 sky130_fd_sc_hd__xor2_1 _17797_ (.A(_01573_),
    .B(_01580_),
    .X(_01581_));
 sky130_fd_sc_hd__xnor2_1 _17798_ (.A(_01567_),
    .B(_01581_),
    .Y(_01582_));
 sky130_fd_sc_hd__xnor2_1 _17799_ (.A(_01566_),
    .B(_01582_),
    .Y(_01583_));
 sky130_fd_sc_hd__nand2_1 _17800_ (.A(_01472_),
    .B(_01474_),
    .Y(_01584_));
 sky130_fd_sc_hd__nor2_1 _17801_ (.A(_09182_),
    .B(_09976_),
    .Y(_01585_));
 sky130_fd_sc_hd__nand2_1 _17802_ (.A(_01472_),
    .B(_01473_),
    .Y(_01586_));
 sky130_fd_sc_hd__mux2_2 _17803_ (.A0(_09182_),
    .A1(_01585_),
    .S(_01586_),
    .X(_01587_));
 sky130_fd_sc_hd__xor2_4 _17804_ (.A(_10111_),
    .B(_01587_),
    .X(_01588_));
 sky130_fd_sc_hd__xor2_1 _17805_ (.A(_01584_),
    .B(_01588_),
    .X(_01589_));
 sky130_fd_sc_hd__xnor2_1 _17806_ (.A(_10121_),
    .B(_01589_),
    .Y(_01590_));
 sky130_fd_sc_hd__inv_2 _17807_ (.A(_10120_),
    .Y(_01591_));
 sky130_fd_sc_hd__nor2_1 _17808_ (.A(_01591_),
    .B(_01480_),
    .Y(_01592_));
 sky130_fd_sc_hd__nor2_1 _17809_ (.A(_01590_),
    .B(_01592_),
    .Y(_01593_));
 sky130_fd_sc_hd__nand2_1 _17810_ (.A(_01590_),
    .B(_01592_),
    .Y(_01594_));
 sky130_fd_sc_hd__and2b_1 _17811_ (.A_N(_01593_),
    .B(_01594_),
    .X(_01595_));
 sky130_fd_sc_hd__xnor2_1 _17812_ (.A(_01583_),
    .B(_01595_),
    .Y(_01596_));
 sky130_fd_sc_hd__a21o_1 _17813_ (.A1(_01470_),
    .A2(_01484_),
    .B1(_01482_),
    .X(_01597_));
 sky130_fd_sc_hd__xnor2_1 _17814_ (.A(_01596_),
    .B(_01597_),
    .Y(_01598_));
 sky130_fd_sc_hd__xnor2_1 _17815_ (.A(_01564_),
    .B(_01598_),
    .Y(_01599_));
 sky130_fd_sc_hd__nor2_1 _17816_ (.A(_01485_),
    .B(_01486_),
    .Y(_01600_));
 sky130_fd_sc_hd__a21oi_1 _17817_ (.A1(_01448_),
    .A2(_01487_),
    .B1(_01600_),
    .Y(_01601_));
 sky130_fd_sc_hd__xor2_1 _17818_ (.A(_01599_),
    .B(_01601_),
    .X(_01602_));
 sky130_fd_sc_hd__xnor2_1 _17819_ (.A(_01524_),
    .B(_01602_),
    .Y(_01603_));
 sky130_fd_sc_hd__a21oi_1 _17820_ (.A1(_10161_),
    .A2(_01493_),
    .B1(_01491_),
    .Y(_01604_));
 sky130_fd_sc_hd__xnor2_1 _17821_ (.A(_01603_),
    .B(_01604_),
    .Y(_01605_));
 sky130_fd_sc_hd__xor2_1 _17822_ (.A(_01515_),
    .B(_01605_),
    .X(_01606_));
 sky130_fd_sc_hd__and3_1 _17823_ (.A(_01513_),
    .B(_01514_),
    .C(_01606_),
    .X(_01607_));
 sky130_fd_sc_hd__a21o_1 _17824_ (.A1(_01513_),
    .A2(_01514_),
    .B1(_01606_),
    .X(_01608_));
 sky130_fd_sc_hd__or2b_2 _17825_ (.A(_01607_),
    .B_N(_01608_),
    .X(_01609_));
 sky130_fd_sc_hd__and3_1 _17826_ (.A(_01498_),
    .B(_01504_),
    .C(_01609_),
    .X(_01610_));
 sky130_fd_sc_hd__a21oi_1 _17827_ (.A1(_01498_),
    .A2(_01504_),
    .B1(_01609_),
    .Y(_01611_));
 sky130_fd_sc_hd__or3_1 _17828_ (.A(_03797_),
    .B(_01610_),
    .C(_01611_),
    .X(_01612_));
 sky130_fd_sc_hd__or2_1 _17829_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .B(\rbzero.wall_tracer.stepDistX[7] ),
    .X(_01613_));
 sky130_fd_sc_hd__nand2_1 _17830_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .B(\rbzero.wall_tracer.stepDistX[7] ),
    .Y(_01614_));
 sky130_fd_sc_hd__o21bai_1 _17831_ (.A1(_01507_),
    .A2(_01509_),
    .B1_N(_01508_),
    .Y(_01615_));
 sky130_fd_sc_hd__a21oi_1 _17832_ (.A1(_01613_),
    .A2(_01614_),
    .B1(_01615_),
    .Y(_01616_));
 sky130_fd_sc_hd__a31o_1 _17833_ (.A1(_01613_),
    .A2(_01614_),
    .A3(_01615_),
    .B1(_09351_),
    .X(_01617_));
 sky130_fd_sc_hd__o21a_1 _17834_ (.A1(_01616_),
    .A2(_01617_),
    .B1(_09275_),
    .X(_01618_));
 sky130_fd_sc_hd__o2bb2a_1 _17835_ (.A1_N(_01612_),
    .A2_N(_01618_),
    .B1(\rbzero.wall_tracer.trackDistX[7] ),
    .B2(_09276_),
    .X(_00560_));
 sky130_fd_sc_hd__a21o_1 _17836_ (.A1(_10121_),
    .A2(_01589_),
    .B1(_01591_),
    .X(_01619_));
 sky130_fd_sc_hd__o21ai_2 _17837_ (.A1(_09182_),
    .A2(_01586_),
    .B1(_01472_),
    .Y(_01620_));
 sky130_fd_sc_hd__xor2_2 _17838_ (.A(_01588_),
    .B(_01620_),
    .X(_01621_));
 sky130_fd_sc_hd__xor2_1 _17839_ (.A(_10121_),
    .B(_01621_),
    .X(_01622_));
 sky130_fd_sc_hd__and2_1 _17840_ (.A(_01619_),
    .B(_01622_),
    .X(_01623_));
 sky130_fd_sc_hd__nor2_1 _17841_ (.A(_01619_),
    .B(_01622_),
    .Y(_01624_));
 sky130_fd_sc_hd__nor2_1 _17842_ (.A(_01623_),
    .B(_01624_),
    .Y(_01625_));
 sky130_fd_sc_hd__nor2_1 _17843_ (.A(_01578_),
    .B(_01579_),
    .Y(_01626_));
 sky130_fd_sc_hd__a21o_1 _17844_ (.A1(_01573_),
    .A2(_01580_),
    .B1(_01626_),
    .X(_01627_));
 sky130_fd_sc_hd__nand2_1 _17845_ (.A(_10111_),
    .B(_01587_),
    .Y(_01628_));
 sky130_fd_sc_hd__a21bo_1 _17846_ (.A1(_01584_),
    .A2(_01588_),
    .B1_N(_01628_),
    .X(_01629_));
 sky130_fd_sc_hd__or4_1 _17847_ (.A(_08594_),
    .B(_09428_),
    .C(_08634_),
    .D(_09462_),
    .X(_01630_));
 sky130_fd_sc_hd__o22ai_1 _17848_ (.A1(_09428_),
    .A2(_08634_),
    .B1(_09463_),
    .B2(_08594_),
    .Y(_01631_));
 sky130_fd_sc_hd__nand2_1 _17849_ (.A(_01630_),
    .B(_01631_),
    .Y(_01632_));
 sky130_fd_sc_hd__or3_1 _17850_ (.A(_07886_),
    .B(_08645_),
    .C(_01632_),
    .X(_01633_));
 sky130_fd_sc_hd__o21ai_1 _17851_ (.A1(_07886_),
    .A2(_08645_),
    .B1(_01632_),
    .Y(_01634_));
 sky130_fd_sc_hd__and2_1 _17852_ (.A(_01633_),
    .B(_01634_),
    .X(_01635_));
 sky130_fd_sc_hd__or2_1 _17853_ (.A(_08240_),
    .B(_09976_),
    .X(_01636_));
 sky130_fd_sc_hd__or2_1 _17854_ (.A(_08241_),
    .B(_01636_),
    .X(_01637_));
 sky130_fd_sc_hd__o2bb2a_1 _17855_ (.A1_N(_01574_),
    .A2_N(_01636_),
    .B1(_01637_),
    .B2(_09978_),
    .X(_01638_));
 sky130_fd_sc_hd__nor2_1 _17856_ (.A(_09968_),
    .B(_09603_),
    .Y(_01639_));
 sky130_fd_sc_hd__xnor2_1 _17857_ (.A(_01638_),
    .B(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hd__o2bb2a_1 _17858_ (.A1_N(_01575_),
    .A2_N(_01577_),
    .B1(_01458_),
    .B2(_01574_),
    .X(_01641_));
 sky130_fd_sc_hd__xor2_1 _17859_ (.A(_01640_),
    .B(_01641_),
    .X(_01642_));
 sky130_fd_sc_hd__xor2_1 _17860_ (.A(_01635_),
    .B(_01642_),
    .X(_01643_));
 sky130_fd_sc_hd__xnor2_1 _17861_ (.A(_01629_),
    .B(_01643_),
    .Y(_01644_));
 sky130_fd_sc_hd__xnor2_2 _17862_ (.A(_01627_),
    .B(_01644_),
    .Y(_01645_));
 sky130_fd_sc_hd__xnor2_2 _17863_ (.A(_01625_),
    .B(_01645_),
    .Y(_01646_));
 sky130_fd_sc_hd__a21oi_2 _17864_ (.A1(_01583_),
    .A2(_01594_),
    .B1(_01593_),
    .Y(_01647_));
 sky130_fd_sc_hd__xor2_2 _17865_ (.A(_01646_),
    .B(_01647_),
    .X(_01648_));
 sky130_fd_sc_hd__a21o_1 _17866_ (.A1(_01547_),
    .A2(_01560_),
    .B1(_01559_),
    .X(_01649_));
 sky130_fd_sc_hd__or2b_1 _17867_ (.A(_01582_),
    .B_N(_01566_),
    .X(_01650_));
 sky130_fd_sc_hd__a21bo_1 _17868_ (.A1(_01567_),
    .A2(_01581_),
    .B1_N(_01650_),
    .X(_01651_));
 sky130_fd_sc_hd__o21ba_1 _17869_ (.A1(_09429_),
    .A2(_08852_),
    .B1_N(_01529_),
    .X(_01652_));
 sky130_fd_sc_hd__or3b_1 _17870_ (.A(_09429_),
    .B(_08851_),
    .C_N(_01529_),
    .X(_01653_));
 sky130_fd_sc_hd__or2b_1 _17871_ (.A(_01652_),
    .B_N(_01653_),
    .X(_01654_));
 sky130_fd_sc_hd__nand2_1 _17872_ (.A(_09684_),
    .B(_09389_),
    .Y(_01655_));
 sky130_fd_sc_hd__xor2_1 _17873_ (.A(_01654_),
    .B(_01655_),
    .X(_01656_));
 sky130_fd_sc_hd__or3_1 _17874_ (.A(_07678_),
    .B(_08531_),
    .C(_01535_),
    .X(_01657_));
 sky130_fd_sc_hd__o21ai_1 _17875_ (.A1(_07678_),
    .A2(_08531_),
    .B1(_01535_),
    .Y(_01658_));
 sky130_fd_sc_hd__nand2_1 _17876_ (.A(_01657_),
    .B(_01658_),
    .Y(_01659_));
 sky130_fd_sc_hd__or2_1 _17877_ (.A(_07670_),
    .B(_08723_),
    .X(_01660_));
 sky130_fd_sc_hd__xnor2_1 _17878_ (.A(_01659_),
    .B(_01660_),
    .Y(_01661_));
 sky130_fd_sc_hd__o31a_1 _17879_ (.A1(_10056_),
    .A2(_08724_),
    .A3(_01534_),
    .B1(_01536_),
    .X(_01662_));
 sky130_fd_sc_hd__or2_1 _17880_ (.A(_01661_),
    .B(_01662_),
    .X(_01663_));
 sky130_fd_sc_hd__nand2_1 _17881_ (.A(_01661_),
    .B(_01662_),
    .Y(_01664_));
 sky130_fd_sc_hd__and2_1 _17882_ (.A(_01663_),
    .B(_01664_),
    .X(_01665_));
 sky130_fd_sc_hd__nand2_1 _17883_ (.A(_01656_),
    .B(_01665_),
    .Y(_01666_));
 sky130_fd_sc_hd__or2_1 _17884_ (.A(_01656_),
    .B(_01665_),
    .X(_01667_));
 sky130_fd_sc_hd__and2_1 _17885_ (.A(_01666_),
    .B(_01667_),
    .X(_01668_));
 sky130_fd_sc_hd__a21bo_1 _17886_ (.A1(_01551_),
    .A2(_01553_),
    .B1_N(_01550_),
    .X(_01669_));
 sky130_fd_sc_hd__nand2_1 _17887_ (.A(_01568_),
    .B(_01571_),
    .Y(_01670_));
 sky130_fd_sc_hd__nor2_1 _17888_ (.A(_07619_),
    .B(_07827_),
    .Y(_01671_));
 sky130_fd_sc_hd__nor2_1 _17889_ (.A(_10095_),
    .B(_08671_),
    .Y(_01672_));
 sky130_fd_sc_hd__xnor2_1 _17890_ (.A(_01671_),
    .B(_01672_),
    .Y(_01673_));
 sky130_fd_sc_hd__or3_1 _17891_ (.A(_09955_),
    .B(_07914_),
    .C(_01673_),
    .X(_01674_));
 sky130_fd_sc_hd__o21ai_1 _17892_ (.A1(_09955_),
    .A2(_07914_),
    .B1(_01673_),
    .Y(_01675_));
 sky130_fd_sc_hd__nand2_1 _17893_ (.A(_01674_),
    .B(_01675_),
    .Y(_01676_));
 sky130_fd_sc_hd__xnor2_1 _17894_ (.A(_01670_),
    .B(_01676_),
    .Y(_01677_));
 sky130_fd_sc_hd__xnor2_1 _17895_ (.A(_01669_),
    .B(_01677_),
    .Y(_01678_));
 sky130_fd_sc_hd__a21oi_1 _17896_ (.A1(_01452_),
    .A2(_01455_),
    .B1(_01554_),
    .Y(_01679_));
 sky130_fd_sc_hd__a21oi_1 _17897_ (.A1(_01548_),
    .A2(_01555_),
    .B1(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__xor2_1 _17898_ (.A(_01678_),
    .B(_01680_),
    .X(_01681_));
 sky130_fd_sc_hd__xnor2_1 _17899_ (.A(_01668_),
    .B(_01681_),
    .Y(_01682_));
 sky130_fd_sc_hd__xor2_1 _17900_ (.A(_01651_),
    .B(_01682_),
    .X(_01683_));
 sky130_fd_sc_hd__xnor2_1 _17901_ (.A(_01649_),
    .B(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__xnor2_1 _17902_ (.A(_01648_),
    .B(_01684_),
    .Y(_01685_));
 sky130_fd_sc_hd__or2b_1 _17903_ (.A(_01596_),
    .B_N(_01597_),
    .X(_01686_));
 sky130_fd_sc_hd__a21boi_2 _17904_ (.A1(_01564_),
    .A2(_01598_),
    .B1_N(_01686_),
    .Y(_01687_));
 sky130_fd_sc_hd__nor2_1 _17905_ (.A(_01685_),
    .B(_01687_),
    .Y(_01688_));
 sky130_fd_sc_hd__and2_1 _17906_ (.A(_01685_),
    .B(_01687_),
    .X(_01689_));
 sky130_fd_sc_hd__nor2_1 _17907_ (.A(_01688_),
    .B(_01689_),
    .Y(_01690_));
 sky130_fd_sc_hd__or2b_1 _17908_ (.A(_01562_),
    .B_N(_01527_),
    .X(_01691_));
 sky130_fd_sc_hd__or2b_1 _17909_ (.A(_01563_),
    .B_N(_01525_),
    .X(_01692_));
 sky130_fd_sc_hd__nand2_1 _17910_ (.A(_01528_),
    .B(_01529_),
    .Y(_01693_));
 sky130_fd_sc_hd__o31a_1 _17911_ (.A1(_08135_),
    .A2(_09115_),
    .A3(_01530_),
    .B1(_01693_),
    .X(_01694_));
 sky130_fd_sc_hd__a21oi_2 _17912_ (.A1(_01542_),
    .A2(_01545_),
    .B1(_01694_),
    .Y(_01695_));
 sky130_fd_sc_hd__and3_1 _17913_ (.A(_01542_),
    .B(_01545_),
    .C(_01694_),
    .X(_01696_));
 sky130_fd_sc_hd__or2_1 _17914_ (.A(_01695_),
    .B(_01696_),
    .X(_01697_));
 sky130_fd_sc_hd__a21o_1 _17915_ (.A1(_01691_),
    .A2(_01692_),
    .B1(_01697_),
    .X(_01698_));
 sky130_fd_sc_hd__nand3_1 _17916_ (.A(_01691_),
    .B(_01692_),
    .C(_01697_),
    .Y(_01699_));
 sky130_fd_sc_hd__and2_1 _17917_ (.A(_01698_),
    .B(_01699_),
    .X(_01700_));
 sky130_fd_sc_hd__xnor2_1 _17918_ (.A(_01518_),
    .B(_01700_),
    .Y(_01701_));
 sky130_fd_sc_hd__xnor2_1 _17919_ (.A(_01690_),
    .B(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__nor2_1 _17920_ (.A(_01599_),
    .B(_01601_),
    .Y(_01703_));
 sky130_fd_sc_hd__a21oi_2 _17921_ (.A1(_01524_),
    .A2(_01602_),
    .B1(_01703_),
    .Y(_01704_));
 sky130_fd_sc_hd__xnor2_1 _17922_ (.A(_01702_),
    .B(_01704_),
    .Y(_01705_));
 sky130_fd_sc_hd__inv_2 _17923_ (.A(_01523_),
    .Y(_01706_));
 sky130_fd_sc_hd__o21a_1 _17924_ (.A1(_10155_),
    .A2(_01706_),
    .B1(_01521_),
    .X(_01707_));
 sky130_fd_sc_hd__xnor2_1 _17925_ (.A(_01705_),
    .B(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hd__or2b_1 _17926_ (.A(_01605_),
    .B_N(_01515_),
    .X(_01709_));
 sky130_fd_sc_hd__o21a_1 _17927_ (.A1(_01603_),
    .A2(_01604_),
    .B1(_01709_),
    .X(_01710_));
 sky130_fd_sc_hd__or2_1 _17928_ (.A(_01708_),
    .B(_01710_),
    .X(_01711_));
 sky130_fd_sc_hd__nand2_1 _17929_ (.A(_01708_),
    .B(_01710_),
    .Y(_01712_));
 sky130_fd_sc_hd__and2_1 _17930_ (.A(_01711_),
    .B(_01712_),
    .X(_01713_));
 sky130_fd_sc_hd__a21oi_2 _17931_ (.A1(_01498_),
    .A2(_01608_),
    .B1(_01607_),
    .Y(_01714_));
 sky130_fd_sc_hd__or2_1 _17932_ (.A(_01502_),
    .B(_01714_),
    .X(_01715_));
 sky130_fd_sc_hd__a31o_2 _17933_ (.A1(_10023_),
    .A2(_10024_),
    .A3(_01501_),
    .B1(_01715_),
    .X(_01716_));
 sky130_fd_sc_hd__o21bai_2 _17934_ (.A1(_01500_),
    .A2(_01609_),
    .B1_N(_01714_),
    .Y(_01717_));
 sky130_fd_sc_hd__and2_1 _17935_ (.A(_01716_),
    .B(_01717_),
    .X(_01718_));
 sky130_fd_sc_hd__nor2_1 _17936_ (.A(_01713_),
    .B(_01718_),
    .Y(_01719_));
 sky130_fd_sc_hd__nand2_1 _17937_ (.A(_01713_),
    .B(_01718_),
    .Y(_01720_));
 sky130_fd_sc_hd__or3b_2 _17938_ (.A(_03797_),
    .B(_01719_),
    .C_N(_01720_),
    .X(_01721_));
 sky130_fd_sc_hd__nor2_1 _17939_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .Y(_01722_));
 sky130_fd_sc_hd__nand2_1 _17940_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .Y(_01723_));
 sky130_fd_sc_hd__and2b_1 _17941_ (.A_N(_01722_),
    .B(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__a21boi_1 _17942_ (.A1(_01613_),
    .A2(_01615_),
    .B1_N(_01614_),
    .Y(_01725_));
 sky130_fd_sc_hd__xnor2_1 _17943_ (.A(_01724_),
    .B(_01725_),
    .Y(_01726_));
 sky130_fd_sc_hd__a21oi_1 _17944_ (.A1(_09279_),
    .A2(_01726_),
    .B1(_09283_),
    .Y(_01727_));
 sky130_fd_sc_hd__o2bb2a_1 _17945_ (.A1_N(_01721_),
    .A2_N(_01727_),
    .B1(\rbzero.wall_tracer.trackDistX[8] ),
    .B2(_09276_),
    .X(_00561_));
 sky130_fd_sc_hd__or2_1 _17946_ (.A(_01702_),
    .B(_01704_),
    .X(_01728_));
 sky130_fd_sc_hd__or2_1 _17947_ (.A(_01705_),
    .B(_01707_),
    .X(_01729_));
 sky130_fd_sc_hd__nor3_2 _17948_ (.A(_09861_),
    .B(_09989_),
    .C(_01621_),
    .Y(_01730_));
 sky130_fd_sc_hd__and2_1 _17949_ (.A(_01591_),
    .B(_01621_),
    .X(_01731_));
 sky130_fd_sc_hd__or2_1 _17950_ (.A(_01730_),
    .B(_01731_),
    .X(_01732_));
 sky130_fd_sc_hd__inv_2 _17951_ (.A(_01732_),
    .Y(_01733_));
 sky130_fd_sc_hd__nor2_1 _17952_ (.A(_01640_),
    .B(_01641_),
    .Y(_01734_));
 sky130_fd_sc_hd__a21o_1 _17953_ (.A1(_01635_),
    .A2(_01642_),
    .B1(_01734_),
    .X(_01735_));
 sky130_fd_sc_hd__a21bo_2 _17954_ (.A1(_01588_),
    .A2(_01620_),
    .B1_N(_01628_),
    .X(_01736_));
 sky130_fd_sc_hd__nor2_1 _17955_ (.A(_08594_),
    .B(_09603_),
    .Y(_01737_));
 sky130_fd_sc_hd__nor2_1 _17956_ (.A(_09428_),
    .B(_08787_),
    .Y(_01738_));
 sky130_fd_sc_hd__xnor2_1 _17957_ (.A(_01737_),
    .B(_01738_),
    .Y(_01739_));
 sky130_fd_sc_hd__or3_1 _17958_ (.A(_07631_),
    .B(_08634_),
    .C(_01739_),
    .X(_01740_));
 sky130_fd_sc_hd__o21ai_1 _17959_ (.A1(_07631_),
    .A2(_08634_),
    .B1(_01739_),
    .Y(_01741_));
 sky130_fd_sc_hd__and2_1 _17960_ (.A(_01740_),
    .B(_01741_),
    .X(_01742_));
 sky130_fd_sc_hd__a21oi_1 _17961_ (.A1(_08240_),
    .A2(_08241_),
    .B1(_09976_),
    .Y(_01743_));
 sky130_fd_sc_hd__nand2_1 _17962_ (.A(_01637_),
    .B(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__nor2_1 _17963_ (.A(_09968_),
    .B(_09978_),
    .Y(_01745_));
 sky130_fd_sc_hd__xor2_1 _17964_ (.A(_01744_),
    .B(_01745_),
    .X(_01746_));
 sky130_fd_sc_hd__o2bb2a_1 _17965_ (.A1_N(_01638_),
    .A2_N(_01639_),
    .B1(_09978_),
    .B2(_01637_),
    .X(_01747_));
 sky130_fd_sc_hd__xor2_1 _17966_ (.A(_01746_),
    .B(_01747_),
    .X(_01748_));
 sky130_fd_sc_hd__nand2_1 _17967_ (.A(_01742_),
    .B(_01748_),
    .Y(_01749_));
 sky130_fd_sc_hd__or2_1 _17968_ (.A(_01742_),
    .B(_01748_),
    .X(_01750_));
 sky130_fd_sc_hd__and2_1 _17969_ (.A(_01749_),
    .B(_01750_),
    .X(_01751_));
 sky130_fd_sc_hd__xnor2_1 _17970_ (.A(_01736_),
    .B(_01751_),
    .Y(_01752_));
 sky130_fd_sc_hd__xnor2_1 _17971_ (.A(_01735_),
    .B(_01752_),
    .Y(_01753_));
 sky130_fd_sc_hd__xnor2_1 _17972_ (.A(_01733_),
    .B(_01753_),
    .Y(_01754_));
 sky130_fd_sc_hd__a21oi_2 _17973_ (.A1(_01625_),
    .A2(_01645_),
    .B1(_01623_),
    .Y(_01755_));
 sky130_fd_sc_hd__xor2_1 _17974_ (.A(_01754_),
    .B(_01755_),
    .X(_01756_));
 sky130_fd_sc_hd__nor2_1 _17975_ (.A(_01678_),
    .B(_01680_),
    .Y(_01757_));
 sky130_fd_sc_hd__a21o_1 _17976_ (.A1(_01668_),
    .A2(_01681_),
    .B1(_01757_),
    .X(_01758_));
 sky130_fd_sc_hd__or2b_1 _17977_ (.A(_01644_),
    .B_N(_01627_),
    .X(_01759_));
 sky130_fd_sc_hd__a21bo_1 _17978_ (.A1(_01629_),
    .A2(_01643_),
    .B1_N(_01759_),
    .X(_01760_));
 sky130_fd_sc_hd__or2_1 _17979_ (.A(_07670_),
    .B(_08851_),
    .X(_01761_));
 sky130_fd_sc_hd__or3_1 _17980_ (.A(_09429_),
    .B(_09373_),
    .C(_01761_),
    .X(_01762_));
 sky130_fd_sc_hd__o21ai_1 _17981_ (.A1(_09429_),
    .A2(_09373_),
    .B1(_01761_),
    .Y(_01763_));
 sky130_fd_sc_hd__nand2_1 _17982_ (.A(_01762_),
    .B(_01763_),
    .Y(_01764_));
 sky130_fd_sc_hd__nor2_1 _17983_ (.A(_08123_),
    .B(_09115_),
    .Y(_01765_));
 sky130_fd_sc_hd__xnor2_1 _17984_ (.A(_01764_),
    .B(_01765_),
    .Y(_01766_));
 sky130_fd_sc_hd__nor2_1 _17985_ (.A(_07678_),
    .B(_08531_),
    .Y(_01767_));
 sky130_fd_sc_hd__nor2_1 _17986_ (.A(_09955_),
    .B(_08663_),
    .Y(_01768_));
 sky130_fd_sc_hd__o22a_1 _17987_ (.A1(_09955_),
    .A2(_08531_),
    .B1(_08985_),
    .B2(_09829_),
    .X(_01769_));
 sky130_fd_sc_hd__a21oi_1 _17988_ (.A1(_01767_),
    .A2(_01768_),
    .B1(_01769_),
    .Y(_01770_));
 sky130_fd_sc_hd__nor2_1 _17989_ (.A(_09833_),
    .B(_08725_),
    .Y(_01771_));
 sky130_fd_sc_hd__xnor2_1 _17990_ (.A(_01770_),
    .B(_01771_),
    .Y(_01772_));
 sky130_fd_sc_hd__o31a_1 _17991_ (.A1(_07760_),
    .A2(_08725_),
    .A3(_01659_),
    .B1(_01657_),
    .X(_01773_));
 sky130_fd_sc_hd__or2_1 _17992_ (.A(_01772_),
    .B(_01773_),
    .X(_01774_));
 sky130_fd_sc_hd__nand2_1 _17993_ (.A(_01772_),
    .B(_01773_),
    .Y(_01775_));
 sky130_fd_sc_hd__and2_1 _17994_ (.A(_01774_),
    .B(_01775_),
    .X(_01776_));
 sky130_fd_sc_hd__nand2_1 _17995_ (.A(_01766_),
    .B(_01776_),
    .Y(_01777_));
 sky130_fd_sc_hd__or2_1 _17996_ (.A(_01766_),
    .B(_01776_),
    .X(_01778_));
 sky130_fd_sc_hd__and2_1 _17997_ (.A(_01777_),
    .B(_01778_),
    .X(_01779_));
 sky130_fd_sc_hd__a21bo_1 _17998_ (.A1(_01671_),
    .A2(_01672_),
    .B1_N(_01674_),
    .X(_01780_));
 sky130_fd_sc_hd__nand2_1 _17999_ (.A(_01630_),
    .B(_01633_),
    .Y(_01781_));
 sky130_fd_sc_hd__nor2_1 _18000_ (.A(_08732_),
    .B(_08645_),
    .Y(_01782_));
 sky130_fd_sc_hd__nor2_1 _18001_ (.A(_07618_),
    .B(_07827_),
    .Y(_01783_));
 sky130_fd_sc_hd__xnor2_1 _18002_ (.A(_01782_),
    .B(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__or3_1 _18003_ (.A(_10095_),
    .B(_08735_),
    .C(_01784_),
    .X(_01785_));
 sky130_fd_sc_hd__o21ai_1 _18004_ (.A1(_10095_),
    .A2(_08735_),
    .B1(_01784_),
    .Y(_01786_));
 sky130_fd_sc_hd__nand2_1 _18005_ (.A(_01785_),
    .B(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__xnor2_1 _18006_ (.A(_01781_),
    .B(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__xnor2_1 _18007_ (.A(_01780_),
    .B(_01788_),
    .Y(_01789_));
 sky130_fd_sc_hd__a21oi_1 _18008_ (.A1(_01568_),
    .A2(_01571_),
    .B1(_01676_),
    .Y(_01790_));
 sky130_fd_sc_hd__a21oi_1 _18009_ (.A1(_01669_),
    .A2(_01677_),
    .B1(_01790_),
    .Y(_01791_));
 sky130_fd_sc_hd__nor2_1 _18010_ (.A(_01789_),
    .B(_01791_),
    .Y(_01792_));
 sky130_fd_sc_hd__and2_1 _18011_ (.A(_01789_),
    .B(_01791_),
    .X(_01793_));
 sky130_fd_sc_hd__nor2_1 _18012_ (.A(_01792_),
    .B(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__xor2_1 _18013_ (.A(_01779_),
    .B(_01794_),
    .X(_01795_));
 sky130_fd_sc_hd__xnor2_1 _18014_ (.A(_01760_),
    .B(_01795_),
    .Y(_01796_));
 sky130_fd_sc_hd__xnor2_1 _18015_ (.A(_01758_),
    .B(_01796_),
    .Y(_01797_));
 sky130_fd_sc_hd__xnor2_1 _18016_ (.A(_01756_),
    .B(_01797_),
    .Y(_01798_));
 sky130_fd_sc_hd__nor2_1 _18017_ (.A(_01646_),
    .B(_01647_),
    .Y(_01799_));
 sky130_fd_sc_hd__a21oi_1 _18018_ (.A1(_01648_),
    .A2(_01684_),
    .B1(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__xor2_1 _18019_ (.A(_01798_),
    .B(_01800_),
    .X(_01801_));
 sky130_fd_sc_hd__or2b_1 _18020_ (.A(_01682_),
    .B_N(_01651_),
    .X(_01802_));
 sky130_fd_sc_hd__or2b_1 _18021_ (.A(_01683_),
    .B_N(_01649_),
    .X(_01803_));
 sky130_fd_sc_hd__o31a_1 _18022_ (.A1(_09018_),
    .A2(_09115_),
    .A3(_01652_),
    .B1(_01653_),
    .X(_01804_));
 sky130_fd_sc_hd__a21o_1 _18023_ (.A1(_01663_),
    .A2(_01666_),
    .B1(_01804_),
    .X(_01805_));
 sky130_fd_sc_hd__nand3_1 _18024_ (.A(_01663_),
    .B(_01666_),
    .C(_01804_),
    .Y(_01806_));
 sky130_fd_sc_hd__nand2_1 _18025_ (.A(_01805_),
    .B(_01806_),
    .Y(_01807_));
 sky130_fd_sc_hd__a21oi_1 _18026_ (.A1(_01802_),
    .A2(_01803_),
    .B1(_01807_),
    .Y(_01808_));
 sky130_fd_sc_hd__and3_1 _18027_ (.A(_01802_),
    .B(_01803_),
    .C(_01807_),
    .X(_01809_));
 sky130_fd_sc_hd__nor2_1 _18028_ (.A(_01808_),
    .B(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__xor2_1 _18029_ (.A(_01695_),
    .B(_01810_),
    .X(_01811_));
 sky130_fd_sc_hd__xnor2_1 _18030_ (.A(_01801_),
    .B(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__a21oi_1 _18031_ (.A1(_01690_),
    .A2(_01701_),
    .B1(_01688_),
    .Y(_01813_));
 sky130_fd_sc_hd__xnor2_1 _18032_ (.A(_01812_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__inv_2 _18033_ (.A(_01700_),
    .Y(_01815_));
 sky130_fd_sc_hd__o21a_1 _18034_ (.A1(_01518_),
    .A2(_01815_),
    .B1(_01698_),
    .X(_01816_));
 sky130_fd_sc_hd__xnor2_1 _18035_ (.A(_01814_),
    .B(_01816_),
    .Y(_01817_));
 sky130_fd_sc_hd__a21oi_1 _18036_ (.A1(_01728_),
    .A2(_01729_),
    .B1(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__and3_1 _18037_ (.A(_01728_),
    .B(_01729_),
    .C(_01817_),
    .X(_01819_));
 sky130_fd_sc_hd__or2_1 _18038_ (.A(_01818_),
    .B(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__a21oi_1 _18039_ (.A1(_01711_),
    .A2(_01720_),
    .B1(_01820_),
    .Y(_01821_));
 sky130_fd_sc_hd__a31o_1 _18040_ (.A1(_01711_),
    .A2(_01720_),
    .A3(_01820_),
    .B1(_03798_),
    .X(_01822_));
 sky130_fd_sc_hd__or2_2 _18041_ (.A(_01821_),
    .B(_01822_),
    .X(_01823_));
 sky130_fd_sc_hd__or2_1 _18042_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .X(_01824_));
 sky130_fd_sc_hd__nand2_1 _18043_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .Y(_01825_));
 sky130_fd_sc_hd__o21ai_1 _18044_ (.A1(_01722_),
    .A2(_01725_),
    .B1(_01723_),
    .Y(_01826_));
 sky130_fd_sc_hd__a21oi_1 _18045_ (.A1(_01824_),
    .A2(_01825_),
    .B1(_01826_),
    .Y(_01827_));
 sky130_fd_sc_hd__a31o_1 _18046_ (.A1(_01824_),
    .A2(_01825_),
    .A3(_01826_),
    .B1(_09351_),
    .X(_01828_));
 sky130_fd_sc_hd__o21a_1 _18047_ (.A1(_01827_),
    .A2(_01828_),
    .B1(_09275_),
    .X(_01829_));
 sky130_fd_sc_hd__o2bb2a_1 _18048_ (.A1_N(_01823_),
    .A2_N(_01829_),
    .B1(\rbzero.wall_tracer.trackDistX[9] ),
    .B2(_09276_),
    .X(_00562_));
 sky130_fd_sc_hd__inv_2 _18049_ (.A(_01820_),
    .Y(_01830_));
 sky130_fd_sc_hd__a21o_1 _18050_ (.A1(_01728_),
    .A2(_01729_),
    .B1(_01817_),
    .X(_01831_));
 sky130_fd_sc_hd__o21a_1 _18051_ (.A1(_01711_),
    .A2(_01819_),
    .B1(_01831_),
    .X(_01832_));
 sky130_fd_sc_hd__inv_2 _18052_ (.A(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__a41o_1 _18053_ (.A1(_01713_),
    .A2(_01716_),
    .A3(_01717_),
    .A4(_01830_),
    .B1(_01833_),
    .X(_01834_));
 sky130_fd_sc_hd__a21o_1 _18054_ (.A1(_01733_),
    .A2(_01753_),
    .B1(_01731_),
    .X(_01835_));
 sky130_fd_sc_hd__or2_1 _18055_ (.A(_01746_),
    .B(_01747_),
    .X(_01836_));
 sky130_fd_sc_hd__nor2_1 _18056_ (.A(_09428_),
    .B(_08923_),
    .Y(_01837_));
 sky130_fd_sc_hd__and3_1 _18057_ (.A(_09163_),
    .B(_09611_),
    .C(_01837_),
    .X(_01838_));
 sky130_fd_sc_hd__a21oi_1 _18058_ (.A1(_09163_),
    .A2(_09611_),
    .B1(_01837_),
    .Y(_01839_));
 sky130_fd_sc_hd__nor2_1 _18059_ (.A(_01838_),
    .B(_01839_),
    .Y(_01840_));
 sky130_fd_sc_hd__nor2_1 _18060_ (.A(_07631_),
    .B(_08787_),
    .Y(_01841_));
 sky130_fd_sc_hd__xnor2_1 _18061_ (.A(_01840_),
    .B(_01841_),
    .Y(_01842_));
 sky130_fd_sc_hd__o31a_1 _18062_ (.A1(_09968_),
    .A2(_09978_),
    .A3(_01744_),
    .B1(_01637_),
    .X(_01843_));
 sky130_fd_sc_hd__nor2_1 _18063_ (.A(_09968_),
    .B(_09976_),
    .Y(_01844_));
 sky130_fd_sc_hd__xnor2_1 _18064_ (.A(_01744_),
    .B(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__xnor2_1 _18065_ (.A(_01843_),
    .B(_01845_),
    .Y(_01846_));
 sky130_fd_sc_hd__xnor2_1 _18066_ (.A(_01842_),
    .B(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__xnor2_1 _18067_ (.A(_01736_),
    .B(_01847_),
    .Y(_01848_));
 sky130_fd_sc_hd__a21oi_1 _18068_ (.A1(_01836_),
    .A2(_01749_),
    .B1(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__and3_1 _18069_ (.A(_01836_),
    .B(_01749_),
    .C(_01848_),
    .X(_01850_));
 sky130_fd_sc_hd__nor2_1 _18070_ (.A(_01849_),
    .B(_01850_),
    .Y(_01851_));
 sky130_fd_sc_hd__xnor2_1 _18071_ (.A(_01732_),
    .B(_01851_),
    .Y(_01852_));
 sky130_fd_sc_hd__xnor2_1 _18072_ (.A(_01835_),
    .B(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__a21o_1 _18073_ (.A1(_01779_),
    .A2(_01794_),
    .B1(_01792_),
    .X(_01854_));
 sky130_fd_sc_hd__or2b_1 _18074_ (.A(_01752_),
    .B_N(_01735_),
    .X(_01855_));
 sky130_fd_sc_hd__a21bo_1 _18075_ (.A1(_01736_),
    .A2(_01751_),
    .B1_N(_01855_),
    .X(_01856_));
 sky130_fd_sc_hd__o22a_1 _18076_ (.A1(_09833_),
    .A2(_08852_),
    .B1(_09373_),
    .B2(_07760_),
    .X(_01857_));
 sky130_fd_sc_hd__or3_1 _18077_ (.A(_09833_),
    .B(_09373_),
    .C(_01761_),
    .X(_01858_));
 sky130_fd_sc_hd__or2b_1 _18078_ (.A(_01857_),
    .B_N(_01858_),
    .X(_01859_));
 sky130_fd_sc_hd__nand2_1 _18079_ (.A(_09429_),
    .B(_09389_),
    .Y(_01860_));
 sky130_fd_sc_hd__xor2_1 _18080_ (.A(_01859_),
    .B(_01860_),
    .X(_01861_));
 sky130_fd_sc_hd__nor2_1 _18081_ (.A(_10095_),
    .B(_08718_),
    .Y(_01862_));
 sky130_fd_sc_hd__xnor2_1 _18082_ (.A(_01768_),
    .B(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__nor2_1 _18083_ (.A(_09829_),
    .B(_08725_),
    .Y(_01864_));
 sky130_fd_sc_hd__xor2_1 _18084_ (.A(_01863_),
    .B(_01864_),
    .X(_01865_));
 sky130_fd_sc_hd__nand2_1 _18085_ (.A(_01767_),
    .B(_01768_),
    .Y(_01866_));
 sky130_fd_sc_hd__o31a_1 _18086_ (.A1(_09833_),
    .A2(_08725_),
    .A3(_01769_),
    .B1(_01866_),
    .X(_01867_));
 sky130_fd_sc_hd__nor2_1 _18087_ (.A(_01865_),
    .B(_01867_),
    .Y(_01868_));
 sky130_fd_sc_hd__and2_1 _18088_ (.A(_01865_),
    .B(_01867_),
    .X(_01869_));
 sky130_fd_sc_hd__nor2_1 _18089_ (.A(_01868_),
    .B(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hd__xnor2_1 _18090_ (.A(_01861_),
    .B(_01870_),
    .Y(_01871_));
 sky130_fd_sc_hd__a21bo_1 _18091_ (.A1(_01782_),
    .A2(_01783_),
    .B1_N(_01785_),
    .X(_01872_));
 sky130_fd_sc_hd__a21bo_1 _18092_ (.A1(_01737_),
    .A2(_01738_),
    .B1_N(_01740_),
    .X(_01873_));
 sky130_fd_sc_hd__nor2_1 _18093_ (.A(_07619_),
    .B(_08634_),
    .Y(_01874_));
 sky130_fd_sc_hd__nor2_1 _18094_ (.A(_08645_),
    .B(_08671_),
    .Y(_01875_));
 sky130_fd_sc_hd__xnor2_1 _18095_ (.A(_01874_),
    .B(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__nor2_1 _18096_ (.A(_07827_),
    .B(_07914_),
    .Y(_01877_));
 sky130_fd_sc_hd__xnor2_1 _18097_ (.A(_01876_),
    .B(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__nand2_1 _18098_ (.A(_01873_),
    .B(_01878_),
    .Y(_01879_));
 sky130_fd_sc_hd__or2_1 _18099_ (.A(_01873_),
    .B(_01878_),
    .X(_01880_));
 sky130_fd_sc_hd__and2_1 _18100_ (.A(_01879_),
    .B(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__xnor2_1 _18101_ (.A(_01872_),
    .B(_01881_),
    .Y(_01882_));
 sky130_fd_sc_hd__a21oi_1 _18102_ (.A1(_01630_),
    .A2(_01633_),
    .B1(_01787_),
    .Y(_01883_));
 sky130_fd_sc_hd__a21oi_1 _18103_ (.A1(_01780_),
    .A2(_01788_),
    .B1(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__xor2_1 _18104_ (.A(_01882_),
    .B(_01884_),
    .X(_01885_));
 sky130_fd_sc_hd__xnor2_1 _18105_ (.A(_01871_),
    .B(_01885_),
    .Y(_01886_));
 sky130_fd_sc_hd__xnor2_1 _18106_ (.A(_01856_),
    .B(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__xnor2_1 _18107_ (.A(_01854_),
    .B(_01887_),
    .Y(_01888_));
 sky130_fd_sc_hd__xor2_1 _18108_ (.A(_01853_),
    .B(_01888_),
    .X(_01889_));
 sky130_fd_sc_hd__nor2_1 _18109_ (.A(_01754_),
    .B(_01755_),
    .Y(_01890_));
 sky130_fd_sc_hd__a21oi_1 _18110_ (.A1(_01756_),
    .A2(_01797_),
    .B1(_01890_),
    .Y(_01891_));
 sky130_fd_sc_hd__xor2_1 _18111_ (.A(_01889_),
    .B(_01891_),
    .X(_01892_));
 sky130_fd_sc_hd__or2b_1 _18112_ (.A(_01796_),
    .B_N(_01758_),
    .X(_01893_));
 sky130_fd_sc_hd__a21bo_1 _18113_ (.A1(_01760_),
    .A2(_01795_),
    .B1_N(_01893_),
    .X(_01894_));
 sky130_fd_sc_hd__o31a_1 _18114_ (.A1(_08123_),
    .A2(_09115_),
    .A3(_01764_),
    .B1(_01762_),
    .X(_01895_));
 sky130_fd_sc_hd__a21o_1 _18115_ (.A1(_01774_),
    .A2(_01777_),
    .B1(_01895_),
    .X(_01896_));
 sky130_fd_sc_hd__nand3_1 _18116_ (.A(_01774_),
    .B(_01777_),
    .C(_01895_),
    .Y(_01897_));
 sky130_fd_sc_hd__and2_1 _18117_ (.A(_01896_),
    .B(_01897_),
    .X(_01898_));
 sky130_fd_sc_hd__xor2_1 _18118_ (.A(_01894_),
    .B(_01898_),
    .X(_01899_));
 sky130_fd_sc_hd__xnor2_1 _18119_ (.A(_01805_),
    .B(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hd__xnor2_1 _18120_ (.A(_01892_),
    .B(_01900_),
    .Y(_01901_));
 sky130_fd_sc_hd__nor2_1 _18121_ (.A(_01798_),
    .B(_01800_),
    .Y(_01902_));
 sky130_fd_sc_hd__a21oi_1 _18122_ (.A1(_01801_),
    .A2(_01811_),
    .B1(_01902_),
    .Y(_01903_));
 sky130_fd_sc_hd__or2_1 _18123_ (.A(_01901_),
    .B(_01903_),
    .X(_01904_));
 sky130_fd_sc_hd__nand2_1 _18124_ (.A(_01901_),
    .B(_01903_),
    .Y(_01905_));
 sky130_fd_sc_hd__nand2_1 _18125_ (.A(_01904_),
    .B(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hd__a21oi_1 _18126_ (.A1(_01695_),
    .A2(_01810_),
    .B1(_01808_),
    .Y(_01907_));
 sky130_fd_sc_hd__xnor2_1 _18127_ (.A(_01906_),
    .B(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__or2_1 _18128_ (.A(_01812_),
    .B(_01813_),
    .X(_01909_));
 sky130_fd_sc_hd__o21a_1 _18129_ (.A1(_01814_),
    .A2(_01816_),
    .B1(_01909_),
    .X(_01910_));
 sky130_fd_sc_hd__nor2_1 _18130_ (.A(_01908_),
    .B(_01910_),
    .Y(_01911_));
 sky130_fd_sc_hd__and2_1 _18131_ (.A(_01908_),
    .B(_01910_),
    .X(_01912_));
 sky130_fd_sc_hd__or2_1 _18132_ (.A(_01911_),
    .B(_01912_),
    .X(_01913_));
 sky130_fd_sc_hd__and2b_1 _18133_ (.A_N(_01834_),
    .B(_01913_),
    .X(_01914_));
 sky130_fd_sc_hd__and2b_1 _18134_ (.A_N(_01913_),
    .B(_01834_),
    .X(_01915_));
 sky130_fd_sc_hd__or3_2 _18135_ (.A(_05121_),
    .B(_01914_),
    .C(_01915_),
    .X(_01916_));
 sky130_fd_sc_hd__nand2_1 _18136_ (.A(_01824_),
    .B(_01826_),
    .Y(_01917_));
 sky130_fd_sc_hd__xnor2_1 _18137_ (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .B(\rbzero.wall_tracer.stepDistX[10] ),
    .Y(_01918_));
 sky130_fd_sc_hd__a21oi_1 _18138_ (.A1(_01825_),
    .A2(_01917_),
    .B1(_01918_),
    .Y(_01919_));
 sky130_fd_sc_hd__a31o_1 _18139_ (.A1(_01825_),
    .A2(_01918_),
    .A3(_01917_),
    .B1(_09351_),
    .X(_01920_));
 sky130_fd_sc_hd__o21a_1 _18140_ (.A1(_01919_),
    .A2(_01920_),
    .B1(_09275_),
    .X(_01921_));
 sky130_fd_sc_hd__o2bb2a_1 _18141_ (.A1_N(_01916_),
    .A2_N(_01921_),
    .B1(\rbzero.wall_tracer.trackDistX[10] ),
    .B2(_09276_),
    .X(_00563_));
 sky130_fd_sc_hd__or2b_1 _18142_ (.A(_01887_),
    .B_N(_01854_),
    .X(_01922_));
 sky130_fd_sc_hd__a21bo_1 _18143_ (.A1(_01856_),
    .A2(_01886_),
    .B1_N(_01922_),
    .X(_01923_));
 sky130_fd_sc_hd__o21a_1 _18144_ (.A1(_01906_),
    .A2(_01907_),
    .B1(_01904_),
    .X(_01924_));
 sky130_fd_sc_hd__a21o_1 _18145_ (.A1(_01861_),
    .A2(_01870_),
    .B1(_01868_),
    .X(_01925_));
 sky130_fd_sc_hd__nor2_1 _18146_ (.A(_08595_),
    .B(_09051_),
    .Y(_01926_));
 sky130_fd_sc_hd__xnor2_1 _18147_ (.A(_01925_),
    .B(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__nor2_1 _18148_ (.A(_08594_),
    .B(_09976_),
    .Y(_01928_));
 sky130_fd_sc_hd__o21a_1 _18149_ (.A1(_01857_),
    .A2(_01860_),
    .B1(_01858_),
    .X(_01929_));
 sky130_fd_sc_hd__xnor2_1 _18150_ (.A(_01928_),
    .B(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__xnor2_1 _18151_ (.A(_01927_),
    .B(_01930_),
    .Y(_01931_));
 sky130_fd_sc_hd__xnor2_1 _18152_ (.A(_01736_),
    .B(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__o21ba_1 _18153_ (.A1(_01730_),
    .A2(_01851_),
    .B1_N(_01731_),
    .X(_01933_));
 sky130_fd_sc_hd__a21oi_1 _18154_ (.A1(_01736_),
    .A2(_01847_),
    .B1(_01849_),
    .Y(_01934_));
 sky130_fd_sc_hd__or2b_1 _18155_ (.A(_01871_),
    .B_N(_01885_),
    .X(_01935_));
 sky130_fd_sc_hd__o21a_1 _18156_ (.A1(_01882_),
    .A2(_01884_),
    .B1(_01935_),
    .X(_01936_));
 sky130_fd_sc_hd__xnor2_1 _18157_ (.A(_01934_),
    .B(_01936_),
    .Y(_01937_));
 sky130_fd_sc_hd__a21bo_1 _18158_ (.A1(_01872_),
    .A2(_01881_),
    .B1_N(_01879_),
    .X(_01938_));
 sky130_fd_sc_hd__a21oi_1 _18159_ (.A1(_01840_),
    .A2(_01841_),
    .B1(_01838_),
    .Y(_01939_));
 sky130_fd_sc_hd__nand2_1 _18160_ (.A(_01874_),
    .B(_01875_),
    .Y(_01940_));
 sky130_fd_sc_hd__o31a_1 _18161_ (.A1(_07827_),
    .A2(_07914_),
    .A3(_01876_),
    .B1(_01940_),
    .X(_01941_));
 sky130_fd_sc_hd__a21o_1 _18162_ (.A1(_08781_),
    .A2(_08784_),
    .B1(_08732_),
    .X(_01942_));
 sky130_fd_sc_hd__nor2_1 _18163_ (.A(_08735_),
    .B(_08645_),
    .Y(_01943_));
 sky130_fd_sc_hd__xor2_1 _18164_ (.A(_01942_),
    .B(_01943_),
    .X(_01944_));
 sky130_fd_sc_hd__xnor2_1 _18165_ (.A(_01941_),
    .B(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__and2b_1 _18166_ (.A_N(_01863_),
    .B(_01864_),
    .X(_01946_));
 sky130_fd_sc_hd__a21oi_1 _18167_ (.A1(_01768_),
    .A2(_01862_),
    .B1(_01946_),
    .Y(_01947_));
 sky130_fd_sc_hd__o22a_1 _18168_ (.A1(_09829_),
    .A2(_08852_),
    .B1(_09373_),
    .B2(_09833_),
    .X(_01948_));
 sky130_fd_sc_hd__or4_1 _18169_ (.A(_09833_),
    .B(_09829_),
    .C(_08852_),
    .D(_09373_),
    .X(_01949_));
 sky130_fd_sc_hd__or2b_1 _18170_ (.A(_01948_),
    .B_N(_01949_),
    .X(_01950_));
 sky130_fd_sc_hd__a21o_1 _18171_ (.A1(_07818_),
    .A2(_07823_),
    .B1(_08718_),
    .X(_01951_));
 sky130_fd_sc_hd__xor2_1 _18172_ (.A(_01950_),
    .B(_01951_),
    .X(_01952_));
 sky130_fd_sc_hd__xnor2_1 _18173_ (.A(_01947_),
    .B(_01952_),
    .Y(_01953_));
 sky130_fd_sc_hd__nand2_1 _18174_ (.A(_07670_),
    .B(_09389_),
    .Y(_01954_));
 sky130_fd_sc_hd__nand2_1 _18175_ (.A(_08536_),
    .B(_08633_),
    .Y(_01955_));
 sky130_fd_sc_hd__xor2_1 _18176_ (.A(_01954_),
    .B(_01955_),
    .X(_01956_));
 sky130_fd_sc_hd__nor2_1 _18177_ (.A(_10095_),
    .B(_08985_),
    .Y(_01957_));
 sky130_fd_sc_hd__nor2_1 _18178_ (.A(_09955_),
    .B(_08725_),
    .Y(_01958_));
 sky130_fd_sc_hd__xnor2_1 _18179_ (.A(_01957_),
    .B(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__xnor2_1 _18180_ (.A(_01956_),
    .B(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hd__xnor2_1 _18181_ (.A(_01953_),
    .B(_01960_),
    .Y(_01961_));
 sky130_fd_sc_hd__xnor2_1 _18182_ (.A(_01945_),
    .B(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__xnor2_1 _18183_ (.A(_01939_),
    .B(_01962_),
    .Y(_01963_));
 sky130_fd_sc_hd__xnor2_1 _18184_ (.A(_01938_),
    .B(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__inv_2 _18185_ (.A(_01846_),
    .Y(_01965_));
 sky130_fd_sc_hd__and2_1 _18186_ (.A(_09968_),
    .B(_01743_),
    .X(_01966_));
 sky130_fd_sc_hd__a311o_1 _18187_ (.A1(_01637_),
    .A2(_01743_),
    .A3(_01745_),
    .B1(_01844_),
    .C1(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__o21a_1 _18188_ (.A1(_01842_),
    .A2(_01965_),
    .B1(_01967_),
    .X(_01968_));
 sky130_fd_sc_hd__a21oi_2 _18189_ (.A1(_08918_),
    .A2(_08921_),
    .B1(_07886_),
    .Y(_01969_));
 sky130_fd_sc_hd__xnor2_1 _18190_ (.A(_01968_),
    .B(_01969_),
    .Y(_01970_));
 sky130_fd_sc_hd__xnor2_1 _18191_ (.A(_01964_),
    .B(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__xnor2_1 _18192_ (.A(_01937_),
    .B(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__xnor2_1 _18193_ (.A(_01933_),
    .B(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__xnor2_1 _18194_ (.A(_01932_),
    .B(_01973_),
    .Y(_01974_));
 sky130_fd_sc_hd__and2b_1 _18195_ (.A_N(_01853_),
    .B(_01888_),
    .X(_01975_));
 sky130_fd_sc_hd__a21o_1 _18196_ (.A1(_01835_),
    .A2(_01852_),
    .B1(_01975_),
    .X(_01976_));
 sky130_fd_sc_hd__nor2_1 _18197_ (.A(_01894_),
    .B(_01898_),
    .Y(_01977_));
 sky130_fd_sc_hd__nand2_1 _18198_ (.A(_01894_),
    .B(_01898_),
    .Y(_01978_));
 sky130_fd_sc_hd__o21a_1 _18199_ (.A1(_01805_),
    .A2(_01977_),
    .B1(_01978_),
    .X(_01979_));
 sky130_fd_sc_hd__xnor2_1 _18200_ (.A(_01976_),
    .B(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__xnor2_1 _18201_ (.A(_01974_),
    .B(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__nor2_1 _18202_ (.A(_01889_),
    .B(_01891_),
    .Y(_01982_));
 sky130_fd_sc_hd__a21oi_1 _18203_ (.A1(_01892_),
    .A2(_01900_),
    .B1(_01982_),
    .Y(_01983_));
 sky130_fd_sc_hd__xnor2_1 _18204_ (.A(_01896_),
    .B(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__xnor2_1 _18205_ (.A(_01981_),
    .B(_01984_),
    .Y(_01985_));
 sky130_fd_sc_hd__xnor2_1 _18206_ (.A(_01924_),
    .B(_01985_),
    .Y(_01986_));
 sky130_fd_sc_hd__xnor2_1 _18207_ (.A(_01923_),
    .B(_01986_),
    .Y(_01987_));
 sky130_fd_sc_hd__o21a_1 _18208_ (.A1(_01911_),
    .A2(_01915_),
    .B1(_01987_),
    .X(_01988_));
 sky130_fd_sc_hd__or3_1 _18209_ (.A(_01911_),
    .B(_01915_),
    .C(_01987_),
    .X(_01989_));
 sky130_fd_sc_hd__or3b_2 _18210_ (.A(_05121_),
    .B(_01988_),
    .C_N(_01989_),
    .X(_01990_));
 sky130_fd_sc_hd__a21o_1 _18211_ (.A1(\rbzero.wall_tracer.trackDistX[10] ),
    .A2(\rbzero.wall_tracer.stepDistX[10] ),
    .B1(_01919_),
    .X(_01991_));
 sky130_fd_sc_hd__xor2_1 _18212_ (.A(\rbzero.wall_tracer.trackDistX[11] ),
    .B(\rbzero.wall_tracer.stepDistX[11] ),
    .X(_01992_));
 sky130_fd_sc_hd__xnor2_1 _18213_ (.A(_01991_),
    .B(_01992_),
    .Y(_01993_));
 sky130_fd_sc_hd__o21a_1 _18214_ (.A1(_07332_),
    .A2(_01993_),
    .B1(_09275_),
    .X(_01994_));
 sky130_fd_sc_hd__o2bb2a_1 _18215_ (.A1_N(_01990_),
    .A2_N(_01994_),
    .B1(\rbzero.wall_tracer.trackDistX[11] ),
    .B2(_09276_),
    .X(_00564_));
 sky130_fd_sc_hd__o21a_4 _18216_ (.A1(_03797_),
    .A2(_08629_),
    .B1(_05027_),
    .X(_01995_));
 sky130_fd_sc_hd__clkbuf_4 _18217_ (.A(_01995_),
    .X(_01996_));
 sky130_fd_sc_hd__clkbuf_4 _18218_ (.A(_05121_),
    .X(_01997_));
 sky130_fd_sc_hd__nand2_1 _18219_ (.A(\rbzero.wall_tracer.trackDistY[-12] ),
    .B(\rbzero.wall_tracer.stepDistY[-12] ),
    .Y(_01998_));
 sky130_fd_sc_hd__or2_1 _18220_ (.A(\rbzero.wall_tracer.trackDistY[-12] ),
    .B(\rbzero.wall_tracer.stepDistY[-12] ),
    .X(_01999_));
 sky130_fd_sc_hd__o21ai_2 _18221_ (.A1(_03797_),
    .A2(_08629_),
    .B1(_05027_),
    .Y(_02000_));
 sky130_fd_sc_hd__clkbuf_4 _18222_ (.A(_02000_),
    .X(_02001_));
 sky130_fd_sc_hd__a31o_1 _18223_ (.A1(_01997_),
    .A2(_01998_),
    .A3(_01999_),
    .B1(_02001_),
    .X(_02002_));
 sky130_fd_sc_hd__o22a_1 _18224_ (.A1(\rbzero.wall_tracer.trackDistY[-12] ),
    .A2(_01996_),
    .B1(_02002_),
    .B2(_09278_),
    .X(_00565_));
 sky130_fd_sc_hd__or2_1 _18225_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .X(_02003_));
 sky130_fd_sc_hd__nand2_1 _18226_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .Y(_02004_));
 sky130_fd_sc_hd__nand3b_1 _18227_ (.A_N(_01998_),
    .B(_02003_),
    .C(_02004_),
    .Y(_02005_));
 sky130_fd_sc_hd__a21bo_1 _18228_ (.A1(_02003_),
    .A2(_02004_),
    .B1_N(_01998_),
    .X(_02006_));
 sky130_fd_sc_hd__a31o_1 _18229_ (.A1(_01997_),
    .A2(_02005_),
    .A3(_02006_),
    .B1(_02001_),
    .X(_02007_));
 sky130_fd_sc_hd__o22a_1 _18230_ (.A1(\rbzero.wall_tracer.trackDistY[-11] ),
    .A2(_01996_),
    .B1(_02007_),
    .B2(_09286_),
    .X(_00566_));
 sky130_fd_sc_hd__and2_1 _18231_ (.A(_02004_),
    .B(_02005_),
    .X(_02008_));
 sky130_fd_sc_hd__nor2_1 _18232_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .Y(_02009_));
 sky130_fd_sc_hd__and2_1 _18233_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .X(_02010_));
 sky130_fd_sc_hd__or3_1 _18234_ (.A(_02008_),
    .B(_02009_),
    .C(_02010_),
    .X(_02011_));
 sky130_fd_sc_hd__o21ai_1 _18235_ (.A1(_02009_),
    .A2(_02010_),
    .B1(_02008_),
    .Y(_02012_));
 sky130_fd_sc_hd__clkbuf_4 _18236_ (.A(_02000_),
    .X(_02013_));
 sky130_fd_sc_hd__a31o_1 _18237_ (.A1(_01997_),
    .A2(_02011_),
    .A3(_02012_),
    .B1(_02013_),
    .X(_02014_));
 sky130_fd_sc_hd__o22a_1 _18238_ (.A1(\rbzero.wall_tracer.trackDistY[-10] ),
    .A2(_01996_),
    .B1(_02014_),
    .B2(_09294_),
    .X(_00567_));
 sky130_fd_sc_hd__or2_1 _18239_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .B(\rbzero.wall_tracer.stepDistY[-9] ),
    .X(_02015_));
 sky130_fd_sc_hd__nand2_1 _18240_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .B(\rbzero.wall_tracer.stepDistY[-9] ),
    .Y(_02016_));
 sky130_fd_sc_hd__o21bai_1 _18241_ (.A1(_02008_),
    .A2(_02009_),
    .B1_N(_02010_),
    .Y(_02017_));
 sky130_fd_sc_hd__nand3_1 _18242_ (.A(_02015_),
    .B(_02016_),
    .C(_02017_),
    .Y(_02018_));
 sky130_fd_sc_hd__a21o_1 _18243_ (.A1(_02015_),
    .A2(_02016_),
    .B1(_02017_),
    .X(_02019_));
 sky130_fd_sc_hd__a31o_1 _18244_ (.A1(_01997_),
    .A2(_02018_),
    .A3(_02019_),
    .B1(_02013_),
    .X(_02020_));
 sky130_fd_sc_hd__o22a_1 _18245_ (.A1(\rbzero.wall_tracer.trackDistY[-9] ),
    .A2(_01996_),
    .B1(_02020_),
    .B2(_09302_),
    .X(_00568_));
 sky130_fd_sc_hd__nor2_1 _18246_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .B(\rbzero.wall_tracer.stepDistY[-8] ),
    .Y(_02021_));
 sky130_fd_sc_hd__and2_1 _18247_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .B(\rbzero.wall_tracer.stepDistY[-8] ),
    .X(_02022_));
 sky130_fd_sc_hd__a21boi_1 _18248_ (.A1(_02015_),
    .A2(_02017_),
    .B1_N(_02016_),
    .Y(_02023_));
 sky130_fd_sc_hd__or3_1 _18249_ (.A(_02021_),
    .B(_02022_),
    .C(_02023_),
    .X(_02024_));
 sky130_fd_sc_hd__o21ai_1 _18250_ (.A1(_02021_),
    .A2(_02022_),
    .B1(_02023_),
    .Y(_02025_));
 sky130_fd_sc_hd__a31o_1 _18251_ (.A1(_01997_),
    .A2(_02024_),
    .A3(_02025_),
    .B1(_02013_),
    .X(_02026_));
 sky130_fd_sc_hd__o22a_1 _18252_ (.A1(\rbzero.wall_tracer.trackDistY[-8] ),
    .A2(_01996_),
    .B1(_02026_),
    .B2(_09310_),
    .X(_00569_));
 sky130_fd_sc_hd__or2_1 _18253_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .B(\rbzero.wall_tracer.stepDistY[-7] ),
    .X(_02027_));
 sky130_fd_sc_hd__nand2_1 _18254_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .B(\rbzero.wall_tracer.stepDistY[-7] ),
    .Y(_02028_));
 sky130_fd_sc_hd__o21bai_1 _18255_ (.A1(_02021_),
    .A2(_02023_),
    .B1_N(_02022_),
    .Y(_02029_));
 sky130_fd_sc_hd__nand3_1 _18256_ (.A(_02027_),
    .B(_02028_),
    .C(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__a21o_1 _18257_ (.A1(_02027_),
    .A2(_02028_),
    .B1(_02029_),
    .X(_02031_));
 sky130_fd_sc_hd__a31o_1 _18258_ (.A1(_01997_),
    .A2(_02030_),
    .A3(_02031_),
    .B1(_02013_),
    .X(_02032_));
 sky130_fd_sc_hd__o22a_1 _18259_ (.A1(\rbzero.wall_tracer.trackDistY[-7] ),
    .A2(_01996_),
    .B1(_02032_),
    .B2(_09317_),
    .X(_00570_));
 sky130_fd_sc_hd__nor2_1 _18260_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .B(\rbzero.wall_tracer.stepDistY[-6] ),
    .Y(_02033_));
 sky130_fd_sc_hd__and2_1 _18261_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .B(\rbzero.wall_tracer.stepDistY[-6] ),
    .X(_02034_));
 sky130_fd_sc_hd__a21boi_1 _18262_ (.A1(_02027_),
    .A2(_02029_),
    .B1_N(_02028_),
    .Y(_02035_));
 sky130_fd_sc_hd__or3_1 _18263_ (.A(_02033_),
    .B(_02034_),
    .C(_02035_),
    .X(_02036_));
 sky130_fd_sc_hd__o21ai_1 _18264_ (.A1(_02033_),
    .A2(_02034_),
    .B1(_02035_),
    .Y(_02037_));
 sky130_fd_sc_hd__a31o_1 _18265_ (.A1(_01997_),
    .A2(_02036_),
    .A3(_02037_),
    .B1(_02013_),
    .X(_02038_));
 sky130_fd_sc_hd__o22a_1 _18266_ (.A1(\rbzero.wall_tracer.trackDistY[-6] ),
    .A2(_01996_),
    .B1(_02038_),
    .B2(_09324_),
    .X(_00571_));
 sky130_fd_sc_hd__clkbuf_4 _18267_ (.A(_01995_),
    .X(_02039_));
 sky130_fd_sc_hd__or2_1 _18268_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .B(\rbzero.wall_tracer.stepDistY[-5] ),
    .X(_02040_));
 sky130_fd_sc_hd__nand2_1 _18269_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .B(\rbzero.wall_tracer.stepDistY[-5] ),
    .Y(_02041_));
 sky130_fd_sc_hd__o21bai_1 _18270_ (.A1(_02033_),
    .A2(_02035_),
    .B1_N(_02034_),
    .Y(_02042_));
 sky130_fd_sc_hd__nand3_1 _18271_ (.A(_02040_),
    .B(_02041_),
    .C(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__a21o_1 _18272_ (.A1(_02040_),
    .A2(_02041_),
    .B1(_02042_),
    .X(_02044_));
 sky130_fd_sc_hd__a31o_1 _18273_ (.A1(_01997_),
    .A2(_02043_),
    .A3(_02044_),
    .B1(_02013_),
    .X(_02045_));
 sky130_fd_sc_hd__o22a_1 _18274_ (.A1(\rbzero.wall_tracer.trackDistY[-5] ),
    .A2(_02039_),
    .B1(_02045_),
    .B2(_09331_),
    .X(_00572_));
 sky130_fd_sc_hd__nor2_1 _18275_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .B(\rbzero.wall_tracer.stepDistY[-4] ),
    .Y(_02046_));
 sky130_fd_sc_hd__nand2_1 _18276_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .B(\rbzero.wall_tracer.stepDistY[-4] ),
    .Y(_02047_));
 sky130_fd_sc_hd__and2b_1 _18277_ (.A_N(_02046_),
    .B(_02047_),
    .X(_02048_));
 sky130_fd_sc_hd__a21boi_1 _18278_ (.A1(_02040_),
    .A2(_02042_),
    .B1_N(_02041_),
    .Y(_02049_));
 sky130_fd_sc_hd__xnor2_1 _18279_ (.A(_02048_),
    .B(_02049_),
    .Y(_02050_));
 sky130_fd_sc_hd__a21o_1 _18280_ (.A1(_09279_),
    .A2(_02050_),
    .B1(_02001_),
    .X(_02051_));
 sky130_fd_sc_hd__o22a_1 _18281_ (.A1(\rbzero.wall_tracer.trackDistY[-4] ),
    .A2(_02039_),
    .B1(_02051_),
    .B2(_09338_),
    .X(_00573_));
 sky130_fd_sc_hd__or2_1 _18282_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .B(\rbzero.wall_tracer.stepDistY[-3] ),
    .X(_02052_));
 sky130_fd_sc_hd__nand2_1 _18283_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .B(\rbzero.wall_tracer.stepDistY[-3] ),
    .Y(_02053_));
 sky130_fd_sc_hd__o21ai_1 _18284_ (.A1(_02046_),
    .A2(_02049_),
    .B1(_02047_),
    .Y(_02054_));
 sky130_fd_sc_hd__and3_1 _18285_ (.A(_02052_),
    .B(_02053_),
    .C(_02054_),
    .X(_02055_));
 sky130_fd_sc_hd__a21oi_1 _18286_ (.A1(_02052_),
    .A2(_02053_),
    .B1(_02054_),
    .Y(_02056_));
 sky130_fd_sc_hd__o311a_1 _18287_ (.A1(_09345_),
    .A2(_02055_),
    .A3(_02056_),
    .B1(_09352_),
    .C1(_01995_),
    .X(_02057_));
 sky130_fd_sc_hd__a21oi_1 _18288_ (.A1(_07275_),
    .A2(_02001_),
    .B1(_02057_),
    .Y(_00574_));
 sky130_fd_sc_hd__nor2_1 _18289_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .Y(_02058_));
 sky130_fd_sc_hd__and2_1 _18290_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .X(_02059_));
 sky130_fd_sc_hd__a21boi_1 _18291_ (.A1(_02052_),
    .A2(_02054_),
    .B1_N(_02053_),
    .Y(_02060_));
 sky130_fd_sc_hd__or3_1 _18292_ (.A(_02058_),
    .B(_02059_),
    .C(_02060_),
    .X(_02061_));
 sky130_fd_sc_hd__o21ai_1 _18293_ (.A1(_02058_),
    .A2(_02059_),
    .B1(_02060_),
    .Y(_02062_));
 sky130_fd_sc_hd__a31o_1 _18294_ (.A1(_01997_),
    .A2(_02061_),
    .A3(_02062_),
    .B1(_02013_),
    .X(_02063_));
 sky130_fd_sc_hd__o22a_1 _18295_ (.A1(\rbzero.wall_tracer.trackDistY[-2] ),
    .A2(_02039_),
    .B1(_02063_),
    .B2(_09354_),
    .X(_00575_));
 sky130_fd_sc_hd__nor2_1 _18296_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .B(\rbzero.wall_tracer.stepDistY[-1] ),
    .Y(_02064_));
 sky130_fd_sc_hd__nor2_1 _18297_ (.A(_04953_),
    .B(_07702_),
    .Y(_02065_));
 sky130_fd_sc_hd__nand2_1 _18298_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .Y(_02066_));
 sky130_fd_sc_hd__o211a_1 _18299_ (.A1(_02064_),
    .A2(_02065_),
    .B1(_02066_),
    .C1(_02061_),
    .X(_02067_));
 sky130_fd_sc_hd__a211oi_2 _18300_ (.A1(_02066_),
    .A2(_02061_),
    .B1(_02064_),
    .C1(_02065_),
    .Y(_02068_));
 sky130_fd_sc_hd__o311a_1 _18301_ (.A1(_09345_),
    .A2(_02067_),
    .A3(_02068_),
    .B1(_09361_),
    .C1(_01995_),
    .X(_02069_));
 sky130_fd_sc_hd__a21oi_1 _18302_ (.A1(_04953_),
    .A2(_02001_),
    .B1(_02069_),
    .Y(_00576_));
 sky130_fd_sc_hd__or2_1 _18303_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .B(\rbzero.wall_tracer.stepDistY[0] ),
    .X(_02070_));
 sky130_fd_sc_hd__nand2_1 _18304_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .B(\rbzero.wall_tracer.stepDistY[0] ),
    .Y(_02071_));
 sky130_fd_sc_hd__o211a_1 _18305_ (.A1(_02065_),
    .A2(_02068_),
    .B1(_02070_),
    .C1(_02071_),
    .X(_02072_));
 sky130_fd_sc_hd__a211oi_1 _18306_ (.A1(_02070_),
    .A2(_02071_),
    .B1(_02065_),
    .C1(_02068_),
    .Y(_02073_));
 sky130_fd_sc_hd__o311a_1 _18307_ (.A1(_09345_),
    .A2(_02072_),
    .A3(_02073_),
    .B1(_09508_),
    .C1(_01995_),
    .X(_02074_));
 sky130_fd_sc_hd__a21oi_1 _18308_ (.A1(_04945_),
    .A2(_02001_),
    .B1(_02074_),
    .Y(_00577_));
 sky130_fd_sc_hd__or2_1 _18309_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .B(\rbzero.wall_tracer.stepDistY[1] ),
    .X(_02075_));
 sky130_fd_sc_hd__nand2_1 _18310_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .B(\rbzero.wall_tracer.stepDistY[1] ),
    .Y(_02076_));
 sky130_fd_sc_hd__a21o_1 _18311_ (.A1(\rbzero.wall_tracer.trackDistY[0] ),
    .A2(\rbzero.wall_tracer.stepDistY[0] ),
    .B1(_02072_),
    .X(_02077_));
 sky130_fd_sc_hd__and3_1 _18312_ (.A(_02075_),
    .B(_02076_),
    .C(_02077_),
    .X(_02078_));
 sky130_fd_sc_hd__inv_2 _18313_ (.A(_02078_),
    .Y(_02079_));
 sky130_fd_sc_hd__a21o_1 _18314_ (.A1(_02075_),
    .A2(_02076_),
    .B1(_02077_),
    .X(_02080_));
 sky130_fd_sc_hd__a31o_1 _18315_ (.A1(_01997_),
    .A2(_02079_),
    .A3(_02080_),
    .B1(_02013_),
    .X(_02081_));
 sky130_fd_sc_hd__o22a_1 _18316_ (.A1(\rbzero.wall_tracer.trackDistY[1] ),
    .A2(_02039_),
    .B1(_02081_),
    .B2(_09641_),
    .X(_00578_));
 sky130_fd_sc_hd__nand2_1 _18317_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .B(\rbzero.wall_tracer.stepDistY[2] ),
    .Y(_02082_));
 sky130_fd_sc_hd__or2_1 _18318_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .B(\rbzero.wall_tracer.stepDistY[2] ),
    .X(_02083_));
 sky130_fd_sc_hd__nand2_1 _18319_ (.A(_02076_),
    .B(_02079_),
    .Y(_02084_));
 sky130_fd_sc_hd__and3_1 _18320_ (.A(_02082_),
    .B(_02083_),
    .C(_02084_),
    .X(_02085_));
 sky130_fd_sc_hd__inv_2 _18321_ (.A(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hd__a21o_1 _18322_ (.A1(_02082_),
    .A2(_02083_),
    .B1(_02084_),
    .X(_02087_));
 sky130_fd_sc_hd__a31o_1 _18323_ (.A1(_05121_),
    .A2(_02086_),
    .A3(_02087_),
    .B1(_02013_),
    .X(_02088_));
 sky130_fd_sc_hd__o22a_1 _18324_ (.A1(\rbzero.wall_tracer.trackDistY[2] ),
    .A2(_02039_),
    .B1(_02088_),
    .B2(_09765_),
    .X(_00579_));
 sky130_fd_sc_hd__nand2_1 _18325_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .B(\rbzero.wall_tracer.stepDistY[3] ),
    .Y(_02089_));
 sky130_fd_sc_hd__or2_1 _18326_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .B(\rbzero.wall_tracer.stepDistY[3] ),
    .X(_02090_));
 sky130_fd_sc_hd__nand2_1 _18327_ (.A(_02082_),
    .B(_02086_),
    .Y(_02091_));
 sky130_fd_sc_hd__a21o_1 _18328_ (.A1(_02089_),
    .A2(_02090_),
    .B1(_02091_),
    .X(_02092_));
 sky130_fd_sc_hd__nand3_1 _18329_ (.A(_02089_),
    .B(_02090_),
    .C(_02091_),
    .Y(_02093_));
 sky130_fd_sc_hd__a31o_1 _18330_ (.A1(_05121_),
    .A2(_02092_),
    .A3(_02093_),
    .B1(_02013_),
    .X(_02094_));
 sky130_fd_sc_hd__o22a_1 _18331_ (.A1(\rbzero.wall_tracer.trackDistY[3] ),
    .A2(_02039_),
    .B1(_02094_),
    .B2(_09888_),
    .X(_00580_));
 sky130_fd_sc_hd__nor2_1 _18332_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .Y(_02095_));
 sky130_fd_sc_hd__and2_1 _18333_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .X(_02096_));
 sky130_fd_sc_hd__a21boi_1 _18334_ (.A1(_02090_),
    .A2(_02091_),
    .B1_N(_02089_),
    .Y(_02097_));
 sky130_fd_sc_hd__nor3_1 _18335_ (.A(_02095_),
    .B(_02096_),
    .C(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__o21a_1 _18336_ (.A1(_02095_),
    .A2(_02096_),
    .B1(_02097_),
    .X(_02099_));
 sky130_fd_sc_hd__o311a_1 _18337_ (.A1(_09351_),
    .A2(_02098_),
    .A3(_02099_),
    .B1(_10028_),
    .C1(_01995_),
    .X(_02100_));
 sky130_fd_sc_hd__a21oi_1 _18338_ (.A1(_05001_),
    .A2(_02001_),
    .B1(_02100_),
    .Y(_00581_));
 sky130_fd_sc_hd__nor2_1 _18339_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .Y(_02101_));
 sky130_fd_sc_hd__and2_1 _18340_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .X(_02102_));
 sky130_fd_sc_hd__o21ba_1 _18341_ (.A1(_02095_),
    .A2(_02097_),
    .B1_N(_02096_),
    .X(_02103_));
 sky130_fd_sc_hd__nor3_1 _18342_ (.A(_02101_),
    .B(_02102_),
    .C(_02103_),
    .Y(_02104_));
 sky130_fd_sc_hd__o21a_1 _18343_ (.A1(_02101_),
    .A2(_02102_),
    .B1(_02103_),
    .X(_02105_));
 sky130_fd_sc_hd__o311a_1 _18344_ (.A1(_09351_),
    .A2(_02104_),
    .A3(_02105_),
    .B1(_10148_),
    .C1(_01995_),
    .X(_02106_));
 sky130_fd_sc_hd__a21oi_1 _18345_ (.A1(_05002_),
    .A2(_02001_),
    .B1(_02106_),
    .Y(_00582_));
 sky130_fd_sc_hd__nor2_1 _18346_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .Y(_02107_));
 sky130_fd_sc_hd__and2_1 _18347_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .X(_02108_));
 sky130_fd_sc_hd__o21ba_1 _18348_ (.A1(_02101_),
    .A2(_02103_),
    .B1_N(_02102_),
    .X(_02109_));
 sky130_fd_sc_hd__or3_1 _18349_ (.A(_02107_),
    .B(_02108_),
    .C(_02109_),
    .X(_02110_));
 sky130_fd_sc_hd__o21ai_1 _18350_ (.A1(_02107_),
    .A2(_02108_),
    .B1(_02109_),
    .Y(_02111_));
 sky130_fd_sc_hd__a31o_1 _18351_ (.A1(_05121_),
    .A2(_02110_),
    .A3(_02111_),
    .B1(_02000_),
    .X(_02112_));
 sky130_fd_sc_hd__o22a_1 _18352_ (.A1(\rbzero.wall_tracer.trackDistY[6] ),
    .A2(_02039_),
    .B1(_02112_),
    .B2(_01506_),
    .X(_00583_));
 sky130_fd_sc_hd__or2_1 _18353_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .X(_02113_));
 sky130_fd_sc_hd__nand2_1 _18354_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .Y(_02114_));
 sky130_fd_sc_hd__o21bai_1 _18355_ (.A1(_02107_),
    .A2(_02109_),
    .B1_N(_02108_),
    .Y(_02115_));
 sky130_fd_sc_hd__a21oi_1 _18356_ (.A1(_02113_),
    .A2(_02114_),
    .B1(_02115_),
    .Y(_02116_));
 sky130_fd_sc_hd__a31o_1 _18357_ (.A1(_02113_),
    .A2(_02114_),
    .A3(_02115_),
    .B1(_04940_),
    .X(_02117_));
 sky130_fd_sc_hd__o211a_1 _18358_ (.A1(_02116_),
    .A2(_02117_),
    .B1(_01612_),
    .C1(_01995_),
    .X(_02118_));
 sky130_fd_sc_hd__a21oi_1 _18359_ (.A1(_04999_),
    .A2(_02001_),
    .B1(_02118_),
    .Y(_00584_));
 sky130_fd_sc_hd__nor2_1 _18360_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .Y(_02119_));
 sky130_fd_sc_hd__nand2_1 _18361_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .Y(_02120_));
 sky130_fd_sc_hd__or2b_1 _18362_ (.A(_02119_),
    .B_N(_02120_),
    .X(_02121_));
 sky130_fd_sc_hd__a21boi_1 _18363_ (.A1(_02113_),
    .A2(_02115_),
    .B1_N(_02114_),
    .Y(_02122_));
 sky130_fd_sc_hd__xnor2_1 _18364_ (.A(_02121_),
    .B(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__o211a_1 _18365_ (.A1(_09345_),
    .A2(_02123_),
    .B1(_01995_),
    .C1(_01721_),
    .X(_02124_));
 sky130_fd_sc_hd__a21oi_1 _18366_ (.A1(_04992_),
    .A2(_02001_),
    .B1(_02124_),
    .Y(_00585_));
 sky130_fd_sc_hd__or2_1 _18367_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .X(_02125_));
 sky130_fd_sc_hd__nand2_1 _18368_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .Y(_02126_));
 sky130_fd_sc_hd__o21ai_1 _18369_ (.A1(_02119_),
    .A2(_02122_),
    .B1(_02120_),
    .Y(_02127_));
 sky130_fd_sc_hd__a21oi_1 _18370_ (.A1(_02125_),
    .A2(_02126_),
    .B1(_02127_),
    .Y(_02128_));
 sky130_fd_sc_hd__a31o_1 _18371_ (.A1(_02125_),
    .A2(_02126_),
    .A3(_02127_),
    .B1(_09351_),
    .X(_02129_));
 sky130_fd_sc_hd__o21a_1 _18372_ (.A1(_02128_),
    .A2(_02129_),
    .B1(_02039_),
    .X(_02130_));
 sky130_fd_sc_hd__o2bb2a_1 _18373_ (.A1_N(_01823_),
    .A2_N(_02130_),
    .B1(_01996_),
    .B2(\rbzero.wall_tracer.trackDistY[9] ),
    .X(_00586_));
 sky130_fd_sc_hd__nand2_1 _18374_ (.A(_02125_),
    .B(_02127_),
    .Y(_02131_));
 sky130_fd_sc_hd__xnor2_1 _18375_ (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .B(\rbzero.wall_tracer.stepDistY[10] ),
    .Y(_02132_));
 sky130_fd_sc_hd__a21oi_1 _18376_ (.A1(_02126_),
    .A2(_02131_),
    .B1(_02132_),
    .Y(_02133_));
 sky130_fd_sc_hd__a31o_1 _18377_ (.A1(_02126_),
    .A2(_02132_),
    .A3(_02131_),
    .B1(_09351_),
    .X(_02134_));
 sky130_fd_sc_hd__o21a_1 _18378_ (.A1(_02133_),
    .A2(_02134_),
    .B1(_02039_),
    .X(_02135_));
 sky130_fd_sc_hd__o2bb2a_1 _18379_ (.A1_N(_01916_),
    .A2_N(_02135_),
    .B1(_01996_),
    .B2(\rbzero.wall_tracer.trackDistY[10] ),
    .X(_00587_));
 sky130_fd_sc_hd__a21o_1 _18380_ (.A1(\rbzero.wall_tracer.trackDistY[10] ),
    .A2(\rbzero.wall_tracer.stepDistY[10] ),
    .B1(_02133_),
    .X(_02136_));
 sky130_fd_sc_hd__xor2_1 _18381_ (.A(\rbzero.wall_tracer.trackDistY[11] ),
    .B(\rbzero.wall_tracer.stepDistY[11] ),
    .X(_02137_));
 sky130_fd_sc_hd__xnor2_1 _18382_ (.A(_02136_),
    .B(_02137_),
    .Y(_02138_));
 sky130_fd_sc_hd__o21a_1 _18383_ (.A1(_07332_),
    .A2(_02138_),
    .B1(_02039_),
    .X(_02139_));
 sky130_fd_sc_hd__o2bb2a_1 _18384_ (.A1_N(_01990_),
    .A2_N(_02139_),
    .B1(_01996_),
    .B2(\rbzero.wall_tracer.trackDistY[11] ),
    .X(_00588_));
 sky130_fd_sc_hd__and4bb_1 _18385_ (.A_N(\rbzero.spi_registers.spi_cmd[1] ),
    .B_N(\rbzero.spi_registers.spi_cmd[3] ),
    .C(\rbzero.spi_registers.spi_cmd[2] ),
    .D(\rbzero.spi_registers.spi_cmd[0] ),
    .X(_02140_));
 sky130_fd_sc_hd__and3_1 _18386_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_03292_),
    .C(_02140_),
    .X(_02141_));
 sky130_fd_sc_hd__mux2_1 _18387_ (.A0(\rbzero.spi_registers.new_vinf ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_02141_),
    .X(_02142_));
 sky130_fd_sc_hd__clkbuf_1 _18388_ (.A(_02142_),
    .X(_00589_));
 sky130_fd_sc_hd__nor2_1 _18389_ (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[-5] ),
    .Y(_02143_));
 sky130_fd_sc_hd__nand2_1 _18390_ (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[-5] ),
    .Y(_02144_));
 sky130_fd_sc_hd__and2b_1 _18391_ (.A_N(_02143_),
    .B(_02144_),
    .X(_02145_));
 sky130_fd_sc_hd__nor2_1 _18392_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[-7] ),
    .Y(_02146_));
 sky130_fd_sc_hd__nand2_1 _18393_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[-8] ),
    .Y(_02147_));
 sky130_fd_sc_hd__nand2_1 _18394_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-9] ),
    .Y(_02148_));
 sky130_fd_sc_hd__or2_1 _18395_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[-8] ),
    .X(_02149_));
 sky130_fd_sc_hd__nand3b_1 _18396_ (.A_N(_02148_),
    .B(_02149_),
    .C(_02147_),
    .Y(_02150_));
 sky130_fd_sc_hd__and2_1 _18397_ (.A(_02147_),
    .B(_02150_),
    .X(_02151_));
 sky130_fd_sc_hd__nand2_1 _18398_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[-7] ),
    .Y(_02152_));
 sky130_fd_sc_hd__o21ai_1 _18399_ (.A1(_02146_),
    .A2(_02151_),
    .B1(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__a21o_1 _18400_ (.A1(\rbzero.debug_overlay.vplaneX[-6] ),
    .A2(\rbzero.wall_tracer.rayAddendX[-6] ),
    .B1(_02153_),
    .X(_02154_));
 sky130_fd_sc_hd__o21ai_1 _18401_ (.A1(\rbzero.debug_overlay.vplaneX[-6] ),
    .A2(\rbzero.wall_tracer.rayAddendX[-6] ),
    .B1(_02154_),
    .Y(_02155_));
 sky130_fd_sc_hd__xnor2_1 _18402_ (.A(_02145_),
    .B(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hd__clkbuf_4 _18403_ (.A(_03729_),
    .X(_02157_));
 sky130_fd_sc_hd__buf_4 _18404_ (.A(_03810_),
    .X(_02158_));
 sky130_fd_sc_hd__a22o_1 _18405_ (.A1(\rbzero.debug_overlay.vplaneX[-9] ),
    .A2(_02157_),
    .B1(_02158_),
    .B2(\rbzero.wall_tracer.rayAddendX[-5] ),
    .X(_02159_));
 sky130_fd_sc_hd__a21o_1 _18406_ (.A1(_09258_),
    .A2(_02156_),
    .B1(_02159_),
    .X(_00590_));
 sky130_fd_sc_hd__nor2_1 _18407_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .Y(_02160_));
 sky130_fd_sc_hd__and2_1 _18408_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .X(_02161_));
 sky130_fd_sc_hd__o21ai_1 _18409_ (.A1(_02143_),
    .A2(_02155_),
    .B1(_02144_),
    .Y(_02162_));
 sky130_fd_sc_hd__or3_1 _18410_ (.A(_02160_),
    .B(_02161_),
    .C(_02162_),
    .X(_02163_));
 sky130_fd_sc_hd__o21ai_1 _18411_ (.A1(_02160_),
    .A2(_02161_),
    .B1(_02162_),
    .Y(_02164_));
 sky130_fd_sc_hd__a21oi_1 _18412_ (.A1(_02163_),
    .A2(_02164_),
    .B1(_02157_),
    .Y(_02165_));
 sky130_fd_sc_hd__clkbuf_4 _18413_ (.A(_09256_),
    .X(_02166_));
 sky130_fd_sc_hd__nand2_1 _18414_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.debug_overlay.vplaneX[-9] ),
    .Y(_02167_));
 sky130_fd_sc_hd__or2_1 _18415_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.debug_overlay.vplaneX[-9] ),
    .X(_02168_));
 sky130_fd_sc_hd__a31o_1 _18416_ (.A1(_02166_),
    .A2(_02167_),
    .A3(_02168_),
    .B1(_09254_),
    .X(_02169_));
 sky130_fd_sc_hd__o22a_1 _18417_ (.A1(\rbzero.wall_tracer.rayAddendX[-4] ),
    .A2(_00013_),
    .B1(_02165_),
    .B2(_02169_),
    .X(_00591_));
 sky130_fd_sc_hd__or2_1 _18418_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_02168_),
    .X(_02170_));
 sky130_fd_sc_hd__nand2_1 _18419_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_02168_),
    .Y(_02171_));
 sky130_fd_sc_hd__nor2_1 _18420_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_02172_));
 sky130_fd_sc_hd__nand2_1 _18421_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_02173_));
 sky130_fd_sc_hd__or2b_1 _18422_ (.A(_02172_),
    .B_N(_02173_),
    .X(_02174_));
 sky130_fd_sc_hd__or2_1 _18423_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .X(_02175_));
 sky130_fd_sc_hd__a21oi_1 _18424_ (.A1(_02175_),
    .A2(_02162_),
    .B1(_02161_),
    .Y(_02176_));
 sky130_fd_sc_hd__xnor2_1 _18425_ (.A(_02174_),
    .B(_02176_),
    .Y(_02177_));
 sky130_fd_sc_hd__nor2_1 _18426_ (.A(_09256_),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__a31o_1 _18427_ (.A1(_09256_),
    .A2(_02170_),
    .A3(_02171_),
    .B1(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__mux2_1 _18428_ (.A0(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A1(_02179_),
    .S(_03812_),
    .X(_02180_));
 sky130_fd_sc_hd__clkbuf_1 _18429_ (.A(_02180_),
    .X(_00592_));
 sky130_fd_sc_hd__or2_1 _18430_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .X(_02181_));
 sky130_fd_sc_hd__nand2_1 _18431_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .Y(_02182_));
 sky130_fd_sc_hd__nand2_1 _18432_ (.A(_02181_),
    .B(_02182_),
    .Y(_02183_));
 sky130_fd_sc_hd__o21ai_1 _18433_ (.A1(_02172_),
    .A2(_02176_),
    .B1(_02173_),
    .Y(_02184_));
 sky130_fd_sc_hd__xor2_1 _18434_ (.A(_02183_),
    .B(_02184_),
    .X(_02185_));
 sky130_fd_sc_hd__nor2_1 _18435_ (.A(_03730_),
    .B(_02185_),
    .Y(_02186_));
 sky130_fd_sc_hd__nand2_1 _18436_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(_02170_),
    .Y(_02187_));
 sky130_fd_sc_hd__or2_1 _18437_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(_02170_),
    .X(_02188_));
 sky130_fd_sc_hd__a31o_1 _18438_ (.A1(_02166_),
    .A2(_02187_),
    .A3(_02188_),
    .B1(_09254_),
    .X(_02189_));
 sky130_fd_sc_hd__o22a_1 _18439_ (.A1(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A2(_00013_),
    .B1(_02186_),
    .B2(_02189_),
    .X(_00593_));
 sky130_fd_sc_hd__or2_1 _18440_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_02190_));
 sky130_fd_sc_hd__buf_2 _18441_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .X(_02191_));
 sky130_fd_sc_hd__nand2_1 _18442_ (.A(_02191_),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_02192_));
 sky130_fd_sc_hd__a21o_1 _18443_ (.A1(\rbzero.debug_overlay.vplaneX[-2] ),
    .A2(\rbzero.wall_tracer.rayAddendX[-2] ),
    .B1(_02184_),
    .X(_02193_));
 sky130_fd_sc_hd__and4_1 _18444_ (.A(_02181_),
    .B(_02190_),
    .C(_02192_),
    .D(_02193_),
    .X(_02194_));
 sky130_fd_sc_hd__inv_2 _18445_ (.A(_02194_),
    .Y(_02195_));
 sky130_fd_sc_hd__a22o_1 _18446_ (.A1(_02190_),
    .A2(_02192_),
    .B1(_02193_),
    .B2(_02181_),
    .X(_02196_));
 sky130_fd_sc_hd__clkbuf_4 _18447_ (.A(_03810_),
    .X(_02197_));
 sky130_fd_sc_hd__or2_1 _18448_ (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .B(\rbzero.debug_overlay.vplaneX[-9] ),
    .X(_02198_));
 sky130_fd_sc_hd__nand2_1 _18449_ (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .B(\rbzero.debug_overlay.vplaneX[-9] ),
    .Y(_02199_));
 sky130_fd_sc_hd__nand2_1 _18450_ (.A(_02198_),
    .B(_02199_),
    .Y(_02200_));
 sky130_fd_sc_hd__xnor2_1 _18451_ (.A(_02188_),
    .B(_02200_),
    .Y(_02201_));
 sky130_fd_sc_hd__a22o_1 _18452_ (.A1(\rbzero.wall_tracer.rayAddendX[-1] ),
    .A2(_02197_),
    .B1(_02201_),
    .B2(_02157_),
    .X(_02202_));
 sky130_fd_sc_hd__a31o_1 _18453_ (.A1(_09261_),
    .A2(_02195_),
    .A3(_02196_),
    .B1(_02202_),
    .X(_00594_));
 sky130_fd_sc_hd__nand2_1 _18454_ (.A(_02192_),
    .B(_02195_),
    .Y(_02203_));
 sky130_fd_sc_hd__or2_1 _18455_ (.A(\rbzero.debug_overlay.vplaneX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_02204_));
 sky130_fd_sc_hd__nand2_1 _18456_ (.A(\rbzero.debug_overlay.vplaneX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_02205_));
 sky130_fd_sc_hd__nand2_1 _18457_ (.A(_02204_),
    .B(_02205_),
    .Y(_02206_));
 sky130_fd_sc_hd__xnor2_1 _18458_ (.A(_02203_),
    .B(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__nand2_1 _18459_ (.A(_02188_),
    .B(_02200_),
    .Y(_02208_));
 sky130_fd_sc_hd__and2_1 _18460_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.debug_overlay.vplaneX[-8] ),
    .X(_02209_));
 sky130_fd_sc_hd__nor2_1 _18461_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.debug_overlay.vplaneX[-8] ),
    .Y(_02210_));
 sky130_fd_sc_hd__o21ai_1 _18462_ (.A1(_02209_),
    .A2(_02210_),
    .B1(_02198_),
    .Y(_02211_));
 sky130_fd_sc_hd__or3_1 _18463_ (.A(_02198_),
    .B(_02209_),
    .C(_02210_),
    .X(_02212_));
 sky130_fd_sc_hd__and2_1 _18464_ (.A(_02211_),
    .B(_02212_),
    .X(_02213_));
 sky130_fd_sc_hd__or2_1 _18465_ (.A(_02208_),
    .B(_02213_),
    .X(_02214_));
 sky130_fd_sc_hd__nand2_1 _18466_ (.A(_02208_),
    .B(_02213_),
    .Y(_02215_));
 sky130_fd_sc_hd__a31o_1 _18467_ (.A1(_03729_),
    .A2(_02214_),
    .A3(_02215_),
    .B1(_02197_),
    .X(_02216_));
 sky130_fd_sc_hd__a21o_1 _18468_ (.A1(_03819_),
    .A2(_02207_),
    .B1(_02216_),
    .X(_02217_));
 sky130_fd_sc_hd__o21a_1 _18469_ (.A1(\rbzero.wall_tracer.rayAddendX[0] ),
    .A2(_00013_),
    .B1(_02217_),
    .X(_00595_));
 sky130_fd_sc_hd__nand2_1 _18470_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_02218_));
 sky130_fd_sc_hd__or2_1 _18471_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_02219_));
 sky130_fd_sc_hd__or2b_1 _18472_ (.A(_02203_),
    .B_N(_02205_),
    .X(_02220_));
 sky130_fd_sc_hd__nand4_2 _18473_ (.A(_02204_),
    .B(_02218_),
    .C(_02219_),
    .D(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__a22o_1 _18474_ (.A1(_02218_),
    .A2(_02219_),
    .B1(_02220_),
    .B2(_02204_),
    .X(_02222_));
 sky130_fd_sc_hd__nor2_1 _18475_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.debug_overlay.vplaneX[-7] ),
    .Y(_02223_));
 sky130_fd_sc_hd__and2_1 _18476_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.debug_overlay.vplaneX[-7] ),
    .X(_02224_));
 sky130_fd_sc_hd__or2_1 _18477_ (.A(_02223_),
    .B(_02224_),
    .X(_02225_));
 sky130_fd_sc_hd__a21o_1 _18478_ (.A1(_02212_),
    .A2(_02215_),
    .B1(_02225_),
    .X(_02226_));
 sky130_fd_sc_hd__nand3_1 _18479_ (.A(_02212_),
    .B(_02215_),
    .C(_02225_),
    .Y(_02227_));
 sky130_fd_sc_hd__nand2_1 _18480_ (.A(_02226_),
    .B(_02227_),
    .Y(_02228_));
 sky130_fd_sc_hd__xnor2_1 _18481_ (.A(_02210_),
    .B(_02228_),
    .Y(_02229_));
 sky130_fd_sc_hd__a22o_1 _18482_ (.A1(\rbzero.wall_tracer.rayAddendX[1] ),
    .A2(_02197_),
    .B1(_02229_),
    .B2(_02157_),
    .X(_02230_));
 sky130_fd_sc_hd__a31o_1 _18483_ (.A1(_09261_),
    .A2(_02221_),
    .A3(_02222_),
    .B1(_02230_),
    .X(_00596_));
 sky130_fd_sc_hd__nand2_1 _18484_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_02231_));
 sky130_fd_sc_hd__or2_1 _18485_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .X(_02232_));
 sky130_fd_sc_hd__nand2_1 _18486_ (.A(_02231_),
    .B(_02232_),
    .Y(_02233_));
 sky130_fd_sc_hd__a21oi_1 _18487_ (.A1(_02218_),
    .A2(_02221_),
    .B1(_02233_),
    .Y(_02234_));
 sky130_fd_sc_hd__a31o_1 _18488_ (.A1(_02218_),
    .A2(_02221_),
    .A3(_02233_),
    .B1(_03729_),
    .X(_02235_));
 sky130_fd_sc_hd__a21bo_1 _18489_ (.A1(_02215_),
    .A2(_02225_),
    .B1_N(_02210_),
    .X(_02236_));
 sky130_fd_sc_hd__and2_1 _18490_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(\rbzero.debug_overlay.vplaneX[-6] ),
    .X(_02237_));
 sky130_fd_sc_hd__nor2_1 _18491_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(\rbzero.debug_overlay.vplaneX[-6] ),
    .Y(_02238_));
 sky130_fd_sc_hd__nor2_1 _18492_ (.A(_02237_),
    .B(_02238_),
    .Y(_02239_));
 sky130_fd_sc_hd__xnor2_1 _18493_ (.A(_02223_),
    .B(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__a21oi_2 _18494_ (.A1(_02226_),
    .A2(_02236_),
    .B1(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__a31o_1 _18495_ (.A1(_02226_),
    .A2(_02240_),
    .A3(_02236_),
    .B1(_03818_),
    .X(_02242_));
 sky130_fd_sc_hd__o21a_1 _18496_ (.A1(_02241_),
    .A2(_02242_),
    .B1(_03811_),
    .X(_02243_));
 sky130_fd_sc_hd__o21ai_1 _18497_ (.A1(_02234_),
    .A2(_02235_),
    .B1(_02243_),
    .Y(_02244_));
 sky130_fd_sc_hd__o21a_1 _18498_ (.A1(\rbzero.wall_tracer.rayAddendX[2] ),
    .A2(_00013_),
    .B1(_02244_),
    .X(_00597_));
 sky130_fd_sc_hd__nand2_1 _18499_ (.A(_02218_),
    .B(_02231_),
    .Y(_02245_));
 sky130_fd_sc_hd__nor2_1 _18500_ (.A(_02221_),
    .B(_02233_),
    .Y(_02246_));
 sky130_fd_sc_hd__buf_2 _18501_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .X(_02247_));
 sky130_fd_sc_hd__nand2_1 _18502_ (.A(_02247_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_02248_));
 sky130_fd_sc_hd__or2_1 _18503_ (.A(_02247_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_02249_));
 sky130_fd_sc_hd__o211ai_2 _18504_ (.A1(_02245_),
    .A2(_02246_),
    .B1(_02248_),
    .C1(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__a211o_1 _18505_ (.A1(_02248_),
    .A2(_02249_),
    .B1(_02245_),
    .C1(_02246_),
    .X(_02251_));
 sky130_fd_sc_hd__xnor2_1 _18506_ (.A(_02191_),
    .B(\rbzero.debug_overlay.vplaneX[-5] ),
    .Y(_02252_));
 sky130_fd_sc_hd__a21oi_1 _18507_ (.A1(_02223_),
    .A2(_02239_),
    .B1(_02241_),
    .Y(_02253_));
 sky130_fd_sc_hd__xnor2_1 _18508_ (.A(_02252_),
    .B(_02253_),
    .Y(_02254_));
 sky130_fd_sc_hd__xnor2_1 _18509_ (.A(_02238_),
    .B(_02254_),
    .Y(_02255_));
 sky130_fd_sc_hd__a22o_1 _18510_ (.A1(\rbzero.wall_tracer.rayAddendX[3] ),
    .A2(_02197_),
    .B1(_02255_),
    .B2(_02157_),
    .X(_02256_));
 sky130_fd_sc_hd__a31o_1 _18511_ (.A1(_09261_),
    .A2(_02250_),
    .A3(_02251_),
    .B1(_02256_),
    .X(_00598_));
 sky130_fd_sc_hd__xnor2_1 _18512_ (.A(_02247_),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .Y(_02257_));
 sky130_fd_sc_hd__a21oi_1 _18513_ (.A1(_02248_),
    .A2(_02250_),
    .B1(_02257_),
    .Y(_02258_));
 sky130_fd_sc_hd__a31o_1 _18514_ (.A1(_02248_),
    .A2(_02250_),
    .A3(_02257_),
    .B1(_09256_),
    .X(_02259_));
 sky130_fd_sc_hd__or2_1 _18515_ (.A(_02252_),
    .B(_02253_),
    .X(_02260_));
 sky130_fd_sc_hd__nor2_1 _18516_ (.A(\rbzero.debug_overlay.vplaneX[0] ),
    .B(\rbzero.debug_overlay.vplaneX[-4] ),
    .Y(_02261_));
 sky130_fd_sc_hd__and2_1 _18517_ (.A(\rbzero.debug_overlay.vplaneX[0] ),
    .B(\rbzero.debug_overlay.vplaneX[-4] ),
    .X(_02262_));
 sky130_fd_sc_hd__o22ai_1 _18518_ (.A1(_02191_),
    .A2(\rbzero.debug_overlay.vplaneX[-5] ),
    .B1(_02261_),
    .B2(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__or4_1 _18519_ (.A(_02191_),
    .B(\rbzero.debug_overlay.vplaneX[-5] ),
    .C(_02261_),
    .D(_02262_),
    .X(_02264_));
 sky130_fd_sc_hd__nand2_1 _18520_ (.A(_02263_),
    .B(_02264_),
    .Y(_02265_));
 sky130_fd_sc_hd__inv_2 _18521_ (.A(_02241_),
    .Y(_02266_));
 sky130_fd_sc_hd__a21bo_1 _18522_ (.A1(_02266_),
    .A2(_02252_),
    .B1_N(_02238_),
    .X(_02267_));
 sky130_fd_sc_hd__and3_1 _18523_ (.A(_02260_),
    .B(_02265_),
    .C(_02267_),
    .X(_02268_));
 sky130_fd_sc_hd__a21o_1 _18524_ (.A1(_02260_),
    .A2(_02267_),
    .B1(_02265_),
    .X(_02269_));
 sky130_fd_sc_hd__nand2_1 _18525_ (.A(_09256_),
    .B(_02269_),
    .Y(_02270_));
 sky130_fd_sc_hd__o22ai_1 _18526_ (.A1(_02258_),
    .A2(_02259_),
    .B1(_02268_),
    .B2(_02270_),
    .Y(_02271_));
 sky130_fd_sc_hd__mux2_1 _18527_ (.A0(\rbzero.wall_tracer.rayAddendX[4] ),
    .A1(_02271_),
    .S(_03812_),
    .X(_02272_));
 sky130_fd_sc_hd__clkbuf_1 _18528_ (.A(_02272_),
    .X(_00599_));
 sky130_fd_sc_hd__or2_1 _18529_ (.A(_02250_),
    .B(_02257_),
    .X(_02273_));
 sky130_fd_sc_hd__buf_2 _18530_ (.A(_02247_),
    .X(_02274_));
 sky130_fd_sc_hd__clkbuf_4 _18531_ (.A(_02274_),
    .X(_02275_));
 sky130_fd_sc_hd__o21ai_1 _18532_ (.A1(\rbzero.wall_tracer.rayAddendX[4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__nand2_1 _18533_ (.A(_02247_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_02277_));
 sky130_fd_sc_hd__or2_1 _18534_ (.A(_02247_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_02278_));
 sky130_fd_sc_hd__nand2_1 _18535_ (.A(_02277_),
    .B(_02278_),
    .Y(_02279_));
 sky130_fd_sc_hd__a21o_1 _18536_ (.A1(_02273_),
    .A2(_02276_),
    .B1(_02279_),
    .X(_02280_));
 sky130_fd_sc_hd__a31oi_1 _18537_ (.A1(_02279_),
    .A2(_02273_),
    .A3(_02276_),
    .B1(_09269_),
    .Y(_02281_));
 sky130_fd_sc_hd__xor2_1 _18538_ (.A(_02247_),
    .B(\rbzero.debug_overlay.vplaneX[-3] ),
    .X(_02282_));
 sky130_fd_sc_hd__xnor2_1 _18539_ (.A(_02261_),
    .B(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__and3_1 _18540_ (.A(_02264_),
    .B(_02269_),
    .C(_02283_),
    .X(_02284_));
 sky130_fd_sc_hd__a21oi_1 _18541_ (.A1(_02264_),
    .A2(_02269_),
    .B1(_02283_),
    .Y(_02285_));
 sky130_fd_sc_hd__nor3_1 _18542_ (.A(_03819_),
    .B(_02284_),
    .C(_02285_),
    .Y(_02286_));
 sky130_fd_sc_hd__a221o_1 _18543_ (.A1(\rbzero.wall_tracer.rayAddendX[5] ),
    .A2(_02158_),
    .B1(_02280_),
    .B2(_02281_),
    .C1(_02286_),
    .X(_00600_));
 sky130_fd_sc_hd__clkbuf_4 _18544_ (.A(_09257_),
    .X(_02287_));
 sky130_fd_sc_hd__xnor2_1 _18545_ (.A(_02247_),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .Y(_02288_));
 sky130_fd_sc_hd__nand3_1 _18546_ (.A(_02277_),
    .B(_02280_),
    .C(_02288_),
    .Y(_02289_));
 sky130_fd_sc_hd__a21o_1 _18547_ (.A1(_02277_),
    .A2(_02280_),
    .B1(_02288_),
    .X(_02290_));
 sky130_fd_sc_hd__nor2_1 _18548_ (.A(_02274_),
    .B(\rbzero.debug_overlay.vplaneX[-2] ),
    .Y(_02291_));
 sky130_fd_sc_hd__and2_1 _18549_ (.A(_02247_),
    .B(\rbzero.debug_overlay.vplaneX[-2] ),
    .X(_02292_));
 sky130_fd_sc_hd__o22ai_1 _18550_ (.A1(_02274_),
    .A2(\rbzero.debug_overlay.vplaneX[-3] ),
    .B1(_02291_),
    .B2(_02292_),
    .Y(_02293_));
 sky130_fd_sc_hd__or3b_1 _18551_ (.A(_02247_),
    .B(\rbzero.debug_overlay.vplaneX[-3] ),
    .C_N(\rbzero.debug_overlay.vplaneX[-2] ),
    .X(_02294_));
 sky130_fd_sc_hd__nand2_1 _18552_ (.A(_02293_),
    .B(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__a21o_1 _18553_ (.A1(_02261_),
    .A2(_02282_),
    .B1(_02285_),
    .X(_02296_));
 sky130_fd_sc_hd__xnor2_1 _18554_ (.A(_02295_),
    .B(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__a22o_1 _18555_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(_02197_),
    .B1(_02297_),
    .B2(_02157_),
    .X(_02298_));
 sky130_fd_sc_hd__a31o_1 _18556_ (.A1(_02287_),
    .A2(_02289_),
    .A3(_02290_),
    .B1(_02298_),
    .X(_00601_));
 sky130_fd_sc_hd__nand2_1 _18557_ (.A(_02274_),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .Y(_02299_));
 sky130_fd_sc_hd__or2_1 _18558_ (.A(_02274_),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_02300_));
 sky130_fd_sc_hd__nor3_1 _18559_ (.A(_02279_),
    .B(_02273_),
    .C(_02288_),
    .Y(_02301_));
 sky130_fd_sc_hd__o41a_1 _18560_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(\rbzero.wall_tracer.rayAddendX[5] ),
    .A3(\rbzero.wall_tracer.rayAddendX[4] ),
    .A4(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_02274_),
    .X(_02302_));
 sky130_fd_sc_hd__a211o_1 _18561_ (.A1(_02299_),
    .A2(_02300_),
    .B1(_02301_),
    .C1(_02302_),
    .X(_02303_));
 sky130_fd_sc_hd__o211ai_2 _18562_ (.A1(_02301_),
    .A2(_02302_),
    .B1(_02299_),
    .C1(_02300_),
    .Y(_02304_));
 sky130_fd_sc_hd__nor2_1 _18563_ (.A(_02274_),
    .B(_02191_),
    .Y(_02305_));
 sky130_fd_sc_hd__and2_1 _18564_ (.A(_02274_),
    .B(_02191_),
    .X(_02306_));
 sky130_fd_sc_hd__o21bai_1 _18565_ (.A1(_02305_),
    .A2(_02306_),
    .B1_N(_02291_),
    .Y(_02307_));
 sky130_fd_sc_hd__nand2_1 _18566_ (.A(_02191_),
    .B(_02291_),
    .Y(_02308_));
 sky130_fd_sc_hd__nand2_1 _18567_ (.A(_02307_),
    .B(_02308_),
    .Y(_02309_));
 sky130_fd_sc_hd__a21boi_1 _18568_ (.A1(_02293_),
    .A2(_02296_),
    .B1_N(_02294_),
    .Y(_02310_));
 sky130_fd_sc_hd__nand2_1 _18569_ (.A(_02309_),
    .B(_02310_),
    .Y(_02311_));
 sky130_fd_sc_hd__or2_1 _18570_ (.A(_02309_),
    .B(_02310_),
    .X(_02312_));
 sky130_fd_sc_hd__a32o_1 _18571_ (.A1(_02166_),
    .A2(_02311_),
    .A3(_02312_),
    .B1(_02158_),
    .B2(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_02313_));
 sky130_fd_sc_hd__a31o_1 _18572_ (.A1(_02287_),
    .A2(_02303_),
    .A3(_02304_),
    .B1(_02313_),
    .X(_00602_));
 sky130_fd_sc_hd__nand2_1 _18573_ (.A(_02275_),
    .B(\rbzero.debug_overlay.vplaneX[0] ),
    .Y(_02314_));
 sky130_fd_sc_hd__or2_1 _18574_ (.A(_02274_),
    .B(\rbzero.debug_overlay.vplaneX[0] ),
    .X(_02315_));
 sky130_fd_sc_hd__a21oi_1 _18575_ (.A1(_02314_),
    .A2(_02315_),
    .B1(_02305_),
    .Y(_02316_));
 sky130_fd_sc_hd__a21o_1 _18576_ (.A1(\rbzero.debug_overlay.vplaneX[0] ),
    .A2(_02305_),
    .B1(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__a21oi_1 _18577_ (.A1(_02308_),
    .A2(_02312_),
    .B1(_02317_),
    .Y(_02318_));
 sky130_fd_sc_hd__a31o_1 _18578_ (.A1(_02308_),
    .A2(_02312_),
    .A3(_02317_),
    .B1(_03818_),
    .X(_02319_));
 sky130_fd_sc_hd__xnor2_1 _18579_ (.A(_02275_),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .Y(_02320_));
 sky130_fd_sc_hd__nand2_1 _18580_ (.A(_02299_),
    .B(_02304_),
    .Y(_02321_));
 sky130_fd_sc_hd__xnor2_1 _18581_ (.A(_02320_),
    .B(_02321_),
    .Y(_02322_));
 sky130_fd_sc_hd__a2bb2o_1 _18582_ (.A1_N(_02318_),
    .A2_N(_02319_),
    .B1(_03818_),
    .B2(_02322_),
    .X(_02323_));
 sky130_fd_sc_hd__mux2_1 _18583_ (.A0(\rbzero.wall_tracer.rayAddendX[8] ),
    .A1(_02323_),
    .S(_03812_),
    .X(_02324_));
 sky130_fd_sc_hd__clkbuf_1 _18584_ (.A(_02324_),
    .X(_00603_));
 sky130_fd_sc_hd__nor2_1 _18585_ (.A(_02304_),
    .B(_02320_),
    .Y(_02325_));
 sky130_fd_sc_hd__o21a_1 _18586_ (.A1(\rbzero.wall_tracer.rayAddendX[8] ),
    .A2(\rbzero.wall_tracer.rayAddendX[7] ),
    .B1(_02275_),
    .X(_02326_));
 sky130_fd_sc_hd__nand2_1 _18587_ (.A(_02275_),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_02327_));
 sky130_fd_sc_hd__or2_1 _18588_ (.A(_02274_),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_02328_));
 sky130_fd_sc_hd__and2_1 _18589_ (.A(_02327_),
    .B(_02328_),
    .X(_02329_));
 sky130_fd_sc_hd__o21ai_1 _18590_ (.A1(_02325_),
    .A2(_02326_),
    .B1(_02329_),
    .Y(_02330_));
 sky130_fd_sc_hd__or3_1 _18591_ (.A(_02329_),
    .B(_02325_),
    .C(_02326_),
    .X(_02331_));
 sky130_fd_sc_hd__and2_1 _18592_ (.A(_02330_),
    .B(_02331_),
    .X(_02332_));
 sky130_fd_sc_hd__a211oi_1 _18593_ (.A1(\rbzero.debug_overlay.vplaneX[0] ),
    .A2(_02191_),
    .B1(_02318_),
    .C1(_02275_),
    .Y(_02333_));
 sky130_fd_sc_hd__a211o_1 _18594_ (.A1(_02315_),
    .A2(_02318_),
    .B1(_02333_),
    .C1(_03818_),
    .X(_02334_));
 sky130_fd_sc_hd__o221a_1 _18595_ (.A1(\rbzero.wall_tracer.rayAddendX[9] ),
    .A2(_03812_),
    .B1(_09269_),
    .B2(_02332_),
    .C1(_02334_),
    .X(_00604_));
 sky130_fd_sc_hd__inv_2 _18596_ (.A(_02275_),
    .Y(_02335_));
 sky130_fd_sc_hd__o211a_1 _18597_ (.A1(_02191_),
    .A2(_02312_),
    .B1(_03729_),
    .C1(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__xnor2_1 _18598_ (.A(_02275_),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_02337_));
 sky130_fd_sc_hd__a21oi_1 _18599_ (.A1(_02327_),
    .A2(_02330_),
    .B1(_02337_),
    .Y(_02338_));
 sky130_fd_sc_hd__a31o_1 _18600_ (.A1(_02327_),
    .A2(_02330_),
    .A3(_02337_),
    .B1(_09269_),
    .X(_02339_));
 sky130_fd_sc_hd__nor2_1 _18601_ (.A(_02338_),
    .B(_02339_),
    .Y(_02340_));
 sky130_fd_sc_hd__a211o_1 _18602_ (.A1(\rbzero.wall_tracer.rayAddendX[10] ),
    .A2(_02158_),
    .B1(_02336_),
    .C1(_02340_),
    .X(_00605_));
 sky130_fd_sc_hd__or3_1 _18603_ (.A(_02335_),
    .B(_05183_),
    .C(_02326_),
    .X(_02341_));
 sky130_fd_sc_hd__and3b_1 _18604_ (.A_N(_02337_),
    .B(_02325_),
    .C(_02329_),
    .X(_02342_));
 sky130_fd_sc_hd__mux2_1 _18605_ (.A0(_02341_),
    .A1(_02275_),
    .S(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__xnor2_1 _18606_ (.A(\rbzero.wall_tracer.rayAddendX[11] ),
    .B(_02343_),
    .Y(_02344_));
 sky130_fd_sc_hd__a221o_1 _18607_ (.A1(\rbzero.wall_tracer.rayAddendX[11] ),
    .A2(_02158_),
    .B1(_09257_),
    .B2(_02344_),
    .C1(_02336_),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _18608_ (.A0(\rbzero.debug_overlay.playerX[0] ),
    .A1(_03742_),
    .S(_03798_),
    .X(_02345_));
 sky130_fd_sc_hd__mux2_1 _18609_ (.A0(\rbzero.map_rom.f4 ),
    .A1(_02345_),
    .S(_09274_),
    .X(_02346_));
 sky130_fd_sc_hd__clkbuf_1 _18610_ (.A(_02346_),
    .X(_00607_));
 sky130_fd_sc_hd__xnor2_1 _18611_ (.A(\rbzero.map_rom.f3 ),
    .B(_07491_),
    .Y(_02347_));
 sky130_fd_sc_hd__or2_1 _18612_ (.A(\rbzero.map_rom.f4 ),
    .B(_02347_),
    .X(_02348_));
 sky130_fd_sc_hd__nand2_1 _18613_ (.A(\rbzero.map_rom.f4 ),
    .B(_02347_),
    .Y(_02349_));
 sky130_fd_sc_hd__and2_1 _18614_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .B(_04940_),
    .X(_02350_));
 sky130_fd_sc_hd__a31o_1 _18615_ (.A1(_03798_),
    .A2(_02348_),
    .A3(_02349_),
    .B1(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__mux2_1 _18616_ (.A0(\rbzero.map_rom.f3 ),
    .A1(_02351_),
    .S(_09274_),
    .X(_02352_));
 sky130_fd_sc_hd__clkbuf_1 _18617_ (.A(_02352_),
    .X(_00608_));
 sky130_fd_sc_hd__xnor2_1 _18618_ (.A(_03736_),
    .B(_07491_),
    .Y(_02353_));
 sky130_fd_sc_hd__o21ai_1 _18619_ (.A1(_03735_),
    .A2(_07491_),
    .B1(_02349_),
    .Y(_02354_));
 sky130_fd_sc_hd__or2_1 _18620_ (.A(_02353_),
    .B(_02354_),
    .X(_02355_));
 sky130_fd_sc_hd__nand2_1 _18621_ (.A(_02353_),
    .B(_02354_),
    .Y(_02356_));
 sky130_fd_sc_hd__and2_1 _18622_ (.A(\rbzero.debug_overlay.playerX[2] ),
    .B(_04940_),
    .X(_02357_));
 sky130_fd_sc_hd__a31o_1 _18623_ (.A1(_03798_),
    .A2(_02355_),
    .A3(_02356_),
    .B1(_02357_),
    .X(_02358_));
 sky130_fd_sc_hd__mux2_1 _18624_ (.A0(_03736_),
    .A1(_02358_),
    .S(_09274_),
    .X(_02359_));
 sky130_fd_sc_hd__clkbuf_1 _18625_ (.A(_02359_),
    .X(_00609_));
 sky130_fd_sc_hd__xnor2_1 _18626_ (.A(\rbzero.map_rom.f1 ),
    .B(_07491_),
    .Y(_02360_));
 sky130_fd_sc_hd__o21a_1 _18627_ (.A1(_03737_),
    .A2(_07491_),
    .B1(_02356_),
    .X(_02361_));
 sky130_fd_sc_hd__xnor2_1 _18628_ (.A(_02360_),
    .B(_02361_),
    .Y(_02362_));
 sky130_fd_sc_hd__mux2_1 _18629_ (.A0(\rbzero.debug_overlay.playerX[3] ),
    .A1(_02362_),
    .S(_03797_),
    .X(_02363_));
 sky130_fd_sc_hd__mux2_1 _18630_ (.A0(\rbzero.map_rom.f1 ),
    .A1(_02363_),
    .S(_09274_),
    .X(_02364_));
 sky130_fd_sc_hd__clkbuf_1 _18631_ (.A(_02364_),
    .X(_00610_));
 sky130_fd_sc_hd__o21a_1 _18632_ (.A1(_03736_),
    .A2(\rbzero.map_rom.f1 ),
    .B1(_02356_),
    .X(_02365_));
 sky130_fd_sc_hd__a21oi_1 _18633_ (.A1(_03746_),
    .A2(_07491_),
    .B1(_02365_),
    .Y(_02366_));
 sky130_fd_sc_hd__o21ai_1 _18634_ (.A1(_07491_),
    .A2(_02356_),
    .B1(_02366_),
    .Y(_02367_));
 sky130_fd_sc_hd__xnor2_1 _18635_ (.A(\rbzero.map_rom.i_col[4] ),
    .B(_02367_),
    .Y(_02368_));
 sky130_fd_sc_hd__mux2_1 _18636_ (.A0(\rbzero.debug_overlay.playerX[4] ),
    .A1(_02368_),
    .S(_03797_),
    .X(_02369_));
 sky130_fd_sc_hd__mux2_1 _18637_ (.A0(\rbzero.map_rom.i_col[4] ),
    .A1(_02369_),
    .S(_09274_),
    .X(_02370_));
 sky130_fd_sc_hd__clkbuf_1 _18638_ (.A(_02370_),
    .X(_00611_));
 sky130_fd_sc_hd__nor2_1 _18639_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .Y(_02371_));
 sky130_fd_sc_hd__and2_1 _18640_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .X(_02372_));
 sky130_fd_sc_hd__nor2_1 _18641_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[-7] ),
    .Y(_02373_));
 sky130_fd_sc_hd__nand2_1 _18642_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[-8] ),
    .Y(_02374_));
 sky130_fd_sc_hd__nand2_1 _18643_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-9] ),
    .Y(_02375_));
 sky130_fd_sc_hd__or2_1 _18644_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[-8] ),
    .X(_02376_));
 sky130_fd_sc_hd__nand3b_1 _18645_ (.A_N(_02375_),
    .B(_02376_),
    .C(_02374_),
    .Y(_02377_));
 sky130_fd_sc_hd__and2_1 _18646_ (.A(_02374_),
    .B(_02377_),
    .X(_02378_));
 sky130_fd_sc_hd__nand2_1 _18647_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[-7] ),
    .Y(_02379_));
 sky130_fd_sc_hd__o21ai_1 _18648_ (.A1(_02373_),
    .A2(_02378_),
    .B1(_02379_),
    .Y(_02380_));
 sky130_fd_sc_hd__a21o_1 _18649_ (.A1(\rbzero.debug_overlay.vplaneY[-6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[-6] ),
    .B1(_02380_),
    .X(_02381_));
 sky130_fd_sc_hd__o21ai_1 _18650_ (.A1(\rbzero.debug_overlay.vplaneY[-6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[-6] ),
    .B1(_02381_),
    .Y(_02382_));
 sky130_fd_sc_hd__or3_1 _18651_ (.A(_02371_),
    .B(_02372_),
    .C(_02382_),
    .X(_02383_));
 sky130_fd_sc_hd__o21ai_1 _18652_ (.A1(_02371_),
    .A2(_02372_),
    .B1(_02382_),
    .Y(_02384_));
 sky130_fd_sc_hd__a22o_1 _18653_ (.A1(\rbzero.debug_overlay.vplaneY[-9] ),
    .A2(_02166_),
    .B1(_02158_),
    .B2(\rbzero.wall_tracer.rayAddendY[-5] ),
    .X(_02385_));
 sky130_fd_sc_hd__a31o_1 _18654_ (.A1(_02287_),
    .A2(_02383_),
    .A3(_02384_),
    .B1(_02385_),
    .X(_00612_));
 sky130_fd_sc_hd__nor2_1 _18655_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .Y(_02386_));
 sky130_fd_sc_hd__and2_1 _18656_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .X(_02387_));
 sky130_fd_sc_hd__nand2_1 _18657_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .Y(_02388_));
 sky130_fd_sc_hd__o21ai_1 _18658_ (.A1(_02371_),
    .A2(_02382_),
    .B1(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__or3_1 _18659_ (.A(_02386_),
    .B(_02387_),
    .C(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__o21ai_1 _18660_ (.A1(_02386_),
    .A2(_02387_),
    .B1(_02389_),
    .Y(_02391_));
 sky130_fd_sc_hd__a21oi_1 _18661_ (.A1(_02390_),
    .A2(_02391_),
    .B1(_02157_),
    .Y(_02392_));
 sky130_fd_sc_hd__or2_1 _18662_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .X(_02393_));
 sky130_fd_sc_hd__nand2_1 _18663_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .Y(_02394_));
 sky130_fd_sc_hd__a31o_1 _18664_ (.A1(_02166_),
    .A2(_02393_),
    .A3(_02394_),
    .B1(_09254_),
    .X(_02395_));
 sky130_fd_sc_hd__o22a_1 _18665_ (.A1(\rbzero.wall_tracer.rayAddendY[-4] ),
    .A2(_00013_),
    .B1(_02392_),
    .B2(_02395_),
    .X(_00613_));
 sky130_fd_sc_hd__or2_1 _18666_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_02393_),
    .X(_02396_));
 sky130_fd_sc_hd__nand2_1 _18667_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_02393_),
    .Y(_02397_));
 sky130_fd_sc_hd__nor2_1 _18668_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_02398_));
 sky130_fd_sc_hd__nand2_1 _18669_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_02399_));
 sky130_fd_sc_hd__or2b_1 _18670_ (.A(_02398_),
    .B_N(_02399_),
    .X(_02400_));
 sky130_fd_sc_hd__or2_1 _18671_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .X(_02401_));
 sky130_fd_sc_hd__a21oi_1 _18672_ (.A1(_02401_),
    .A2(_02389_),
    .B1(_02387_),
    .Y(_02402_));
 sky130_fd_sc_hd__xnor2_1 _18673_ (.A(_02400_),
    .B(_02402_),
    .Y(_02403_));
 sky130_fd_sc_hd__nor2_1 _18674_ (.A(_09256_),
    .B(_02403_),
    .Y(_02404_));
 sky130_fd_sc_hd__a31o_1 _18675_ (.A1(_09256_),
    .A2(_02396_),
    .A3(_02397_),
    .B1(_02404_),
    .X(_02405_));
 sky130_fd_sc_hd__mux2_1 _18676_ (.A0(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A1(_02405_),
    .S(_03812_),
    .X(_02406_));
 sky130_fd_sc_hd__clkbuf_1 _18677_ (.A(_02406_),
    .X(_00614_));
 sky130_fd_sc_hd__or2_1 _18678_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .X(_02407_));
 sky130_fd_sc_hd__nand2_1 _18679_ (.A(_04260_),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .Y(_02408_));
 sky130_fd_sc_hd__nand2_1 _18680_ (.A(_02407_),
    .B(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__o21ai_1 _18681_ (.A1(_02398_),
    .A2(_02402_),
    .B1(_02399_),
    .Y(_02410_));
 sky130_fd_sc_hd__xor2_1 _18682_ (.A(_02409_),
    .B(_02410_),
    .X(_02411_));
 sky130_fd_sc_hd__nor2_1 _18683_ (.A(_02157_),
    .B(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__nand2_1 _18684_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(_02396_),
    .Y(_02413_));
 sky130_fd_sc_hd__or2_1 _18685_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(_02396_),
    .X(_02414_));
 sky130_fd_sc_hd__a31o_1 _18686_ (.A1(_02166_),
    .A2(_02413_),
    .A3(_02414_),
    .B1(_09254_),
    .X(_02415_));
 sky130_fd_sc_hd__o22a_1 _18687_ (.A1(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A2(_00013_),
    .B1(_02412_),
    .B2(_02415_),
    .X(_00615_));
 sky130_fd_sc_hd__or2_1 _18688_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_02416_));
 sky130_fd_sc_hd__nand2_1 _18689_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_02417_));
 sky130_fd_sc_hd__a21o_1 _18690_ (.A1(_04260_),
    .A2(\rbzero.wall_tracer.rayAddendY[-2] ),
    .B1(_02410_),
    .X(_02418_));
 sky130_fd_sc_hd__and4_1 _18691_ (.A(_02407_),
    .B(_02416_),
    .C(_02417_),
    .D(_02418_),
    .X(_02419_));
 sky130_fd_sc_hd__inv_2 _18692_ (.A(_02419_),
    .Y(_02420_));
 sky130_fd_sc_hd__a22o_1 _18693_ (.A1(_02416_),
    .A2(_02417_),
    .B1(_02418_),
    .B2(_02407_),
    .X(_02421_));
 sky130_fd_sc_hd__or2_1 _18694_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .X(_02422_));
 sky130_fd_sc_hd__nand2_1 _18695_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .Y(_02423_));
 sky130_fd_sc_hd__nand2_1 _18696_ (.A(_02422_),
    .B(_02423_),
    .Y(_02424_));
 sky130_fd_sc_hd__xnor2_1 _18697_ (.A(_02414_),
    .B(_02424_),
    .Y(_02425_));
 sky130_fd_sc_hd__a22o_1 _18698_ (.A1(\rbzero.wall_tracer.rayAddendY[-1] ),
    .A2(_02197_),
    .B1(_02425_),
    .B2(_02157_),
    .X(_02426_));
 sky130_fd_sc_hd__a31o_1 _18699_ (.A1(_02287_),
    .A2(_02420_),
    .A3(_02421_),
    .B1(_02426_),
    .X(_00616_));
 sky130_fd_sc_hd__nand2_1 _18700_ (.A(_02417_),
    .B(_02420_),
    .Y(_02427_));
 sky130_fd_sc_hd__buf_2 _18701_ (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .X(_02428_));
 sky130_fd_sc_hd__nor2_1 _18702_ (.A(_02428_),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .Y(_02429_));
 sky130_fd_sc_hd__and2_1 _18703_ (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_02430_));
 sky130_fd_sc_hd__nor2_1 _18704_ (.A(_02429_),
    .B(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__o21ai_1 _18705_ (.A1(_02427_),
    .A2(_02431_),
    .B1(_03818_),
    .Y(_02432_));
 sky130_fd_sc_hd__a21oi_1 _18706_ (.A1(_02427_),
    .A2(_02431_),
    .B1(_02432_),
    .Y(_02433_));
 sky130_fd_sc_hd__nand2_1 _18707_ (.A(_02414_),
    .B(_02424_),
    .Y(_02434_));
 sky130_fd_sc_hd__and2_1 _18708_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .X(_02435_));
 sky130_fd_sc_hd__nor2_1 _18709_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .Y(_02436_));
 sky130_fd_sc_hd__nor2_1 _18710_ (.A(_02435_),
    .B(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__xnor2_1 _18711_ (.A(_02422_),
    .B(_02437_),
    .Y(_02438_));
 sky130_fd_sc_hd__or2_1 _18712_ (.A(_02434_),
    .B(_02438_),
    .X(_02439_));
 sky130_fd_sc_hd__nand2_1 _18713_ (.A(_02434_),
    .B(_02438_),
    .Y(_02440_));
 sky130_fd_sc_hd__a31o_1 _18714_ (.A1(_02166_),
    .A2(_02439_),
    .A3(_02440_),
    .B1(_09254_),
    .X(_02441_));
 sky130_fd_sc_hd__o22a_1 _18715_ (.A1(\rbzero.wall_tracer.rayAddendY[0] ),
    .A2(_00013_),
    .B1(_02433_),
    .B2(_02441_),
    .X(_00617_));
 sky130_fd_sc_hd__or2_1 _18716_ (.A(_02428_),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_02442_));
 sky130_fd_sc_hd__nand2_1 _18717_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .Y(_02443_));
 sky130_fd_sc_hd__or2_1 _18718_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_02444_));
 sky130_fd_sc_hd__or2_1 _18719_ (.A(_02427_),
    .B(_02430_),
    .X(_02445_));
 sky130_fd_sc_hd__nand4_2 _18720_ (.A(_02442_),
    .B(_02443_),
    .C(_02444_),
    .D(_02445_),
    .Y(_02446_));
 sky130_fd_sc_hd__a22o_1 _18721_ (.A1(_02443_),
    .A2(_02444_),
    .B1(_02445_),
    .B2(_02442_),
    .X(_02447_));
 sky130_fd_sc_hd__or2_1 _18722_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.debug_overlay.vplaneY[-7] ),
    .X(_02448_));
 sky130_fd_sc_hd__nand2_1 _18723_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.debug_overlay.vplaneY[-7] ),
    .Y(_02449_));
 sky130_fd_sc_hd__nand2_1 _18724_ (.A(_02448_),
    .B(_02449_),
    .Y(_02450_));
 sky130_fd_sc_hd__o31ai_1 _18725_ (.A1(_02422_),
    .A2(_02435_),
    .A3(_02436_),
    .B1(_02440_),
    .Y(_02451_));
 sky130_fd_sc_hd__xor2_1 _18726_ (.A(_02450_),
    .B(_02451_),
    .X(_02452_));
 sky130_fd_sc_hd__xnor2_1 _18727_ (.A(_02436_),
    .B(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__a22o_1 _18728_ (.A1(\rbzero.wall_tracer.rayAddendY[1] ),
    .A2(_02197_),
    .B1(_02453_),
    .B2(_02157_),
    .X(_02454_));
 sky130_fd_sc_hd__a31o_1 _18729_ (.A1(_02287_),
    .A2(_02446_),
    .A3(_02447_),
    .B1(_02454_),
    .X(_00618_));
 sky130_fd_sc_hd__nand2_1 _18730_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_02455_));
 sky130_fd_sc_hd__or2_1 _18731_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .X(_02456_));
 sky130_fd_sc_hd__nand2_1 _18732_ (.A(_02455_),
    .B(_02456_),
    .Y(_02457_));
 sky130_fd_sc_hd__a21oi_1 _18733_ (.A1(_02443_),
    .A2(_02446_),
    .B1(_02457_),
    .Y(_02458_));
 sky130_fd_sc_hd__a31o_1 _18734_ (.A1(_02443_),
    .A2(_02446_),
    .A3(_02457_),
    .B1(_09256_),
    .X(_02459_));
 sky130_fd_sc_hd__nand2_1 _18735_ (.A(_04260_),
    .B(\rbzero.debug_overlay.vplaneY[-6] ),
    .Y(_02460_));
 sky130_fd_sc_hd__or2_1 _18736_ (.A(_04260_),
    .B(\rbzero.debug_overlay.vplaneY[-6] ),
    .X(_02461_));
 sky130_fd_sc_hd__nor2_1 _18737_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.debug_overlay.vplaneY[-7] ),
    .Y(_02462_));
 sky130_fd_sc_hd__a21oi_1 _18738_ (.A1(_02460_),
    .A2(_02461_),
    .B1(_02462_),
    .Y(_02463_));
 sky130_fd_sc_hd__and3_1 _18739_ (.A(_02462_),
    .B(_02460_),
    .C(_02461_),
    .X(_02464_));
 sky130_fd_sc_hd__nor2_1 _18740_ (.A(_02463_),
    .B(_02464_),
    .Y(_02465_));
 sky130_fd_sc_hd__nand2_1 _18741_ (.A(_02440_),
    .B(_02450_),
    .Y(_02466_));
 sky130_fd_sc_hd__a32o_1 _18742_ (.A1(_02448_),
    .A2(_02449_),
    .A3(_02451_),
    .B1(_02466_),
    .B2(_02436_),
    .X(_02467_));
 sky130_fd_sc_hd__and2_1 _18743_ (.A(_02465_),
    .B(_02467_),
    .X(_02468_));
 sky130_fd_sc_hd__o21ai_1 _18744_ (.A1(_02465_),
    .A2(_02467_),
    .B1(_09256_),
    .Y(_02469_));
 sky130_fd_sc_hd__o22ai_1 _18745_ (.A1(_02458_),
    .A2(_02459_),
    .B1(_02468_),
    .B2(_02469_),
    .Y(_02470_));
 sky130_fd_sc_hd__mux2_1 _18746_ (.A0(\rbzero.wall_tracer.rayAddendY[2] ),
    .A1(_02470_),
    .S(_03811_),
    .X(_02471_));
 sky130_fd_sc_hd__clkbuf_1 _18747_ (.A(_02471_),
    .X(_00619_));
 sky130_fd_sc_hd__buf_2 _18748_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .X(_02472_));
 sky130_fd_sc_hd__nand2_1 _18749_ (.A(_02472_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_02473_));
 sky130_fd_sc_hd__or2_1 _18750_ (.A(_02472_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_02474_));
 sky130_fd_sc_hd__nand2_1 _18751_ (.A(_02443_),
    .B(_02455_),
    .Y(_02475_));
 sky130_fd_sc_hd__nor2_1 _18752_ (.A(_02446_),
    .B(_02457_),
    .Y(_02476_));
 sky130_fd_sc_hd__a211o_1 _18753_ (.A1(_02473_),
    .A2(_02474_),
    .B1(_02475_),
    .C1(_02476_),
    .X(_02477_));
 sky130_fd_sc_hd__o211ai_2 _18754_ (.A1(_02475_),
    .A2(_02476_),
    .B1(_02473_),
    .C1(_02474_),
    .Y(_02478_));
 sky130_fd_sc_hd__nor2_1 _18755_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.debug_overlay.vplaneY[-5] ),
    .Y(_02479_));
 sky130_fd_sc_hd__and2_1 _18756_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.debug_overlay.vplaneY[-5] ),
    .X(_02480_));
 sky130_fd_sc_hd__nor2_1 _18757_ (.A(_02479_),
    .B(_02480_),
    .Y(_02481_));
 sky130_fd_sc_hd__o21a_1 _18758_ (.A1(_02464_),
    .A2(_02468_),
    .B1(_02481_),
    .X(_02482_));
 sky130_fd_sc_hd__nor3_1 _18759_ (.A(_02464_),
    .B(_02468_),
    .C(_02481_),
    .Y(_02483_));
 sky130_fd_sc_hd__or3_1 _18760_ (.A(_02461_),
    .B(_02482_),
    .C(_02483_),
    .X(_02484_));
 sky130_fd_sc_hd__o21ai_1 _18761_ (.A1(_02482_),
    .A2(_02483_),
    .B1(_02461_),
    .Y(_02485_));
 sky130_fd_sc_hd__a32o_1 _18762_ (.A1(_02166_),
    .A2(_02484_),
    .A3(_02485_),
    .B1(_02158_),
    .B2(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_02486_));
 sky130_fd_sc_hd__a31o_1 _18763_ (.A1(_02287_),
    .A2(_02477_),
    .A3(_02478_),
    .B1(_02486_),
    .X(_00620_));
 sky130_fd_sc_hd__xnor2_1 _18764_ (.A(_02472_),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_02487_));
 sky130_fd_sc_hd__a21oi_1 _18765_ (.A1(_02473_),
    .A2(_02478_),
    .B1(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__a31o_1 _18766_ (.A1(_02473_),
    .A2(_02478_),
    .A3(_02487_),
    .B1(_03729_),
    .X(_02489_));
 sky130_fd_sc_hd__nor2_1 _18767_ (.A(_02488_),
    .B(_02489_),
    .Y(_02490_));
 sky130_fd_sc_hd__xor2_1 _18768_ (.A(_02428_),
    .B(\rbzero.debug_overlay.vplaneY[-4] ),
    .X(_02491_));
 sky130_fd_sc_hd__xor2_1 _18769_ (.A(_02479_),
    .B(_02491_),
    .X(_02492_));
 sky130_fd_sc_hd__nor2_1 _18770_ (.A(_04260_),
    .B(\rbzero.debug_overlay.vplaneY[-6] ),
    .Y(_02493_));
 sky130_fd_sc_hd__o22a_1 _18771_ (.A1(_02468_),
    .A2(_02481_),
    .B1(_02482_),
    .B2(_02493_),
    .X(_02494_));
 sky130_fd_sc_hd__and2_1 _18772_ (.A(_02492_),
    .B(_02494_),
    .X(_02495_));
 sky130_fd_sc_hd__o21ai_1 _18773_ (.A1(_02492_),
    .A2(_02494_),
    .B1(_02166_),
    .Y(_02496_));
 sky130_fd_sc_hd__o21ai_1 _18774_ (.A1(_02495_),
    .A2(_02496_),
    .B1(_03812_),
    .Y(_02497_));
 sky130_fd_sc_hd__o22a_1 _18775_ (.A1(\rbzero.wall_tracer.rayAddendY[4] ),
    .A2(_03812_),
    .B1(_02490_),
    .B2(_02497_),
    .X(_00621_));
 sky130_fd_sc_hd__nor2_1 _18776_ (.A(_02472_),
    .B(\rbzero.debug_overlay.vplaneY[-3] ),
    .Y(_02498_));
 sky130_fd_sc_hd__and2_1 _18777_ (.A(_02472_),
    .B(\rbzero.debug_overlay.vplaneY[-3] ),
    .X(_02499_));
 sky130_fd_sc_hd__o22a_1 _18778_ (.A1(_02428_),
    .A2(\rbzero.debug_overlay.vplaneY[-4] ),
    .B1(_02498_),
    .B2(_02499_),
    .X(_02500_));
 sky130_fd_sc_hd__nor4_1 _18779_ (.A(_02428_),
    .B(\rbzero.debug_overlay.vplaneY[-4] ),
    .C(_02498_),
    .D(_02499_),
    .Y(_02501_));
 sky130_fd_sc_hd__nor2_1 _18780_ (.A(_02500_),
    .B(_02501_),
    .Y(_02502_));
 sky130_fd_sc_hd__a21oi_1 _18781_ (.A1(_02479_),
    .A2(_02491_),
    .B1(_02495_),
    .Y(_02503_));
 sky130_fd_sc_hd__xnor2_1 _18782_ (.A(_02502_),
    .B(_02503_),
    .Y(_02504_));
 sky130_fd_sc_hd__nand2_1 _18783_ (.A(_02472_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_02505_));
 sky130_fd_sc_hd__or2_1 _18784_ (.A(_02472_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_02506_));
 sky130_fd_sc_hd__nand2_1 _18785_ (.A(_02505_),
    .B(_02506_),
    .Y(_02507_));
 sky130_fd_sc_hd__or2_1 _18786_ (.A(_02478_),
    .B(_02487_),
    .X(_02508_));
 sky130_fd_sc_hd__buf_2 _18787_ (.A(_02472_),
    .X(_02509_));
 sky130_fd_sc_hd__buf_2 _18788_ (.A(_02509_),
    .X(_02510_));
 sky130_fd_sc_hd__o21ai_1 _18789_ (.A1(\rbzero.wall_tracer.rayAddendY[4] ),
    .A2(\rbzero.wall_tracer.rayAddendY[3] ),
    .B1(_02510_),
    .Y(_02511_));
 sky130_fd_sc_hd__nand3_1 _18790_ (.A(_02507_),
    .B(_02508_),
    .C(_02511_),
    .Y(_02512_));
 sky130_fd_sc_hd__a21o_1 _18791_ (.A1(_02508_),
    .A2(_02511_),
    .B1(_02507_),
    .X(_02513_));
 sky130_fd_sc_hd__and3_1 _18792_ (.A(_03818_),
    .B(_02512_),
    .C(_02513_),
    .X(_02514_));
 sky130_fd_sc_hd__a21o_1 _18793_ (.A1(_03729_),
    .A2(_02504_),
    .B1(_02514_),
    .X(_02515_));
 sky130_fd_sc_hd__mux2_1 _18794_ (.A0(\rbzero.wall_tracer.rayAddendY[5] ),
    .A1(_02515_),
    .S(_03811_),
    .X(_02516_));
 sky130_fd_sc_hd__clkbuf_1 _18795_ (.A(_02516_),
    .X(_00622_));
 sky130_fd_sc_hd__xnor2_1 _18796_ (.A(_02472_),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_02517_));
 sky130_fd_sc_hd__nand3_1 _18797_ (.A(_02505_),
    .B(_02513_),
    .C(_02517_),
    .Y(_02518_));
 sky130_fd_sc_hd__a21o_1 _18798_ (.A1(_02505_),
    .A2(_02513_),
    .B1(_02517_),
    .X(_02519_));
 sky130_fd_sc_hd__or2_1 _18799_ (.A(_02472_),
    .B(_04260_),
    .X(_02520_));
 sky130_fd_sc_hd__nand2_1 _18800_ (.A(_02509_),
    .B(_04260_),
    .Y(_02521_));
 sky130_fd_sc_hd__a21o_1 _18801_ (.A1(_02520_),
    .A2(_02521_),
    .B1(_02498_),
    .X(_02522_));
 sky130_fd_sc_hd__nand2_1 _18802_ (.A(_04260_),
    .B(_02498_),
    .Y(_02523_));
 sky130_fd_sc_hd__nand2_1 _18803_ (.A(_02522_),
    .B(_02523_),
    .Y(_02524_));
 sky130_fd_sc_hd__o21bai_1 _18804_ (.A1(_02500_),
    .A2(_02503_),
    .B1_N(_02501_),
    .Y(_02525_));
 sky130_fd_sc_hd__xnor2_1 _18805_ (.A(_02524_),
    .B(_02525_),
    .Y(_02526_));
 sky130_fd_sc_hd__a22o_1 _18806_ (.A1(\rbzero.wall_tracer.rayAddendY[6] ),
    .A2(_02197_),
    .B1(_02526_),
    .B2(_02166_),
    .X(_02527_));
 sky130_fd_sc_hd__a31o_1 _18807_ (.A1(_02287_),
    .A2(_02518_),
    .A3(_02519_),
    .B1(_02527_),
    .X(_00623_));
 sky130_fd_sc_hd__nand2_1 _18808_ (.A(_02509_),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .Y(_02528_));
 sky130_fd_sc_hd__or2_1 _18809_ (.A(_02509_),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_02529_));
 sky130_fd_sc_hd__nor3_1 _18810_ (.A(_02507_),
    .B(_02508_),
    .C(_02517_),
    .Y(_02530_));
 sky130_fd_sc_hd__o41a_1 _18811_ (.A1(\rbzero.wall_tracer.rayAddendY[6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[5] ),
    .A3(\rbzero.wall_tracer.rayAddendY[4] ),
    .A4(\rbzero.wall_tracer.rayAddendY[3] ),
    .B1(_02509_),
    .X(_02531_));
 sky130_fd_sc_hd__a211o_1 _18812_ (.A1(_02528_),
    .A2(_02529_),
    .B1(_02530_),
    .C1(_02531_),
    .X(_02532_));
 sky130_fd_sc_hd__o211ai_1 _18813_ (.A1(_02530_),
    .A2(_02531_),
    .B1(_02528_),
    .C1(_02529_),
    .Y(_02533_));
 sky130_fd_sc_hd__or2b_1 _18814_ (.A(_02524_),
    .B_N(_02525_),
    .X(_02534_));
 sky130_fd_sc_hd__nor2_1 _18815_ (.A(_02509_),
    .B(\rbzero.debug_overlay.vplaneY[-1] ),
    .Y(_02535_));
 sky130_fd_sc_hd__and2_1 _18816_ (.A(_02509_),
    .B(\rbzero.debug_overlay.vplaneY[-1] ),
    .X(_02536_));
 sky130_fd_sc_hd__o21ai_1 _18817_ (.A1(_02535_),
    .A2(_02536_),
    .B1(_02520_),
    .Y(_02537_));
 sky130_fd_sc_hd__or3_1 _18818_ (.A(_02520_),
    .B(_02535_),
    .C(_02536_),
    .X(_02538_));
 sky130_fd_sc_hd__nand2_1 _18819_ (.A(_02537_),
    .B(_02538_),
    .Y(_02539_));
 sky130_fd_sc_hd__nand3_1 _18820_ (.A(_02523_),
    .B(_02534_),
    .C(_02539_),
    .Y(_02540_));
 sky130_fd_sc_hd__a21o_1 _18821_ (.A1(_02523_),
    .A2(_02534_),
    .B1(_02539_),
    .X(_02541_));
 sky130_fd_sc_hd__a31o_1 _18822_ (.A1(_03729_),
    .A2(_02540_),
    .A3(_02541_),
    .B1(_02197_),
    .X(_02542_));
 sky130_fd_sc_hd__a31o_1 _18823_ (.A1(_03819_),
    .A2(_02532_),
    .A3(_02533_),
    .B1(_02542_),
    .X(_02543_));
 sky130_fd_sc_hd__o21a_1 _18824_ (.A1(\rbzero.wall_tracer.rayAddendY[7] ),
    .A2(_00013_),
    .B1(_02543_),
    .X(_00624_));
 sky130_fd_sc_hd__xor2_1 _18825_ (.A(_02509_),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .X(_02544_));
 sky130_fd_sc_hd__nand2_1 _18826_ (.A(_02528_),
    .B(_02533_),
    .Y(_02545_));
 sky130_fd_sc_hd__xnor2_1 _18827_ (.A(_02544_),
    .B(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__nand2_1 _18828_ (.A(_02510_),
    .B(_02428_),
    .Y(_02547_));
 sky130_fd_sc_hd__or2_1 _18829_ (.A(_02509_),
    .B(_02428_),
    .X(_02548_));
 sky130_fd_sc_hd__a21oi_1 _18830_ (.A1(_02547_),
    .A2(_02548_),
    .B1(_02535_),
    .Y(_02549_));
 sky130_fd_sc_hd__a21o_1 _18831_ (.A1(_02428_),
    .A2(_02535_),
    .B1(_02549_),
    .X(_02550_));
 sky130_fd_sc_hd__and3_1 _18832_ (.A(_02538_),
    .B(_02541_),
    .C(_02550_),
    .X(_02551_));
 sky130_fd_sc_hd__a21oi_1 _18833_ (.A1(_02538_),
    .A2(_02541_),
    .B1(_02550_),
    .Y(_02552_));
 sky130_fd_sc_hd__or3_1 _18834_ (.A(_03818_),
    .B(_02551_),
    .C(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__o211a_1 _18835_ (.A1(_03729_),
    .A2(_02546_),
    .B1(_02553_),
    .C1(_03812_),
    .X(_02554_));
 sky130_fd_sc_hd__o21ba_1 _18836_ (.A1(\rbzero.wall_tracer.rayAddendY[8] ),
    .A2(_00013_),
    .B1_N(_02554_),
    .X(_00625_));
 sky130_fd_sc_hd__and2b_1 _18837_ (.A_N(_02533_),
    .B(_02544_),
    .X(_02555_));
 sky130_fd_sc_hd__o21a_1 _18838_ (.A1(\rbzero.wall_tracer.rayAddendY[8] ),
    .A2(\rbzero.wall_tracer.rayAddendY[7] ),
    .B1(_02509_),
    .X(_02556_));
 sky130_fd_sc_hd__xor2_1 _18839_ (.A(_02510_),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .X(_02557_));
 sky130_fd_sc_hd__o21a_1 _18840_ (.A1(_02555_),
    .A2(_02556_),
    .B1(_02557_),
    .X(_02558_));
 sky130_fd_sc_hd__nor3_1 _18841_ (.A(_02557_),
    .B(_02555_),
    .C(_02556_),
    .Y(_02559_));
 sky130_fd_sc_hd__nor2_1 _18842_ (.A(_02558_),
    .B(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__a211oi_1 _18843_ (.A1(_02428_),
    .A2(\rbzero.debug_overlay.vplaneY[-1] ),
    .B1(_02552_),
    .C1(_02510_),
    .Y(_02561_));
 sky130_fd_sc_hd__a211o_1 _18844_ (.A1(_02548_),
    .A2(_02552_),
    .B1(_02561_),
    .C1(_03818_),
    .X(_02562_));
 sky130_fd_sc_hd__o221a_1 _18845_ (.A1(\rbzero.wall_tracer.rayAddendY[9] ),
    .A2(_03812_),
    .B1(_09269_),
    .B2(_02560_),
    .C1(_02562_),
    .X(_00626_));
 sky130_fd_sc_hd__a21o_1 _18846_ (.A1(_02510_),
    .A2(\rbzero.wall_tracer.rayAddendY[9] ),
    .B1(_02558_),
    .X(_02563_));
 sky130_fd_sc_hd__xor2_1 _18847_ (.A(_02510_),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .X(_02564_));
 sky130_fd_sc_hd__nand2_1 _18848_ (.A(_02563_),
    .B(_02564_),
    .Y(_02565_));
 sky130_fd_sc_hd__or2_1 _18849_ (.A(_02563_),
    .B(_02564_),
    .X(_02566_));
 sky130_fd_sc_hd__nor2_1 _18850_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_02541_),
    .Y(_02567_));
 sky130_fd_sc_hd__or3_1 _18851_ (.A(_02510_),
    .B(_03818_),
    .C(_02567_),
    .X(_02568_));
 sky130_fd_sc_hd__a21bo_1 _18852_ (.A1(\rbzero.wall_tracer.rayAddendY[10] ),
    .A2(_02158_),
    .B1_N(_02568_),
    .X(_02569_));
 sky130_fd_sc_hd__a31o_1 _18853_ (.A1(_02287_),
    .A2(_02565_),
    .A3(_02566_),
    .B1(_02569_),
    .X(_00627_));
 sky130_fd_sc_hd__or4b_1 _18854_ (.A(\rbzero.wall_tracer.rayAddendY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .C(_02556_),
    .D_N(_02510_),
    .X(_02570_));
 sky130_fd_sc_hd__and3_1 _18855_ (.A(_02557_),
    .B(_02555_),
    .C(_02564_),
    .X(_02571_));
 sky130_fd_sc_hd__mux2_1 _18856_ (.A0(_02570_),
    .A1(_02510_),
    .S(_02571_),
    .X(_02572_));
 sky130_fd_sc_hd__nor2_1 _18857_ (.A(_03809_),
    .B(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__xnor2_1 _18858_ (.A(\rbzero.wall_tracer.rayAddendY[11] ),
    .B(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__o21ai_1 _18859_ (.A1(_03730_),
    .A2(_02574_),
    .B1(_02568_),
    .Y(_00628_));
 sky130_fd_sc_hd__and2b_1 _18860_ (.A_N(\rbzero.spi_registers.sclk_buffer[2] ),
    .B(\rbzero.spi_registers.sclk_buffer[1] ),
    .X(_02575_));
 sky130_fd_sc_hd__clkbuf_2 _18861_ (.A(_02575_),
    .X(_02576_));
 sky130_fd_sc_hd__or3_1 _18862_ (.A(\rbzero.spi_registers.spi_counter[6] ),
    .B(\rbzero.spi_registers.spi_counter[5] ),
    .C(\rbzero.spi_registers.spi_counter[4] ),
    .X(_02577_));
 sky130_fd_sc_hd__or2_1 _18863_ (.A(\rbzero.spi_registers.spi_cmd[1] ),
    .B(\rbzero.spi_registers.spi_cmd[0] ),
    .X(_02578_));
 sky130_fd_sc_hd__a21o_1 _18864_ (.A1(\rbzero.spi_registers.spi_cmd[2] ),
    .A2(_02578_),
    .B1(\rbzero.spi_registers.spi_cmd[3] ),
    .X(_02579_));
 sky130_fd_sc_hd__mux2_1 _18865_ (.A0(\rbzero.spi_registers.spi_counter[3] ),
    .A1(_02579_),
    .S(\rbzero.spi_registers.spi_counter[0] ),
    .X(_02580_));
 sky130_fd_sc_hd__inv_2 _18866_ (.A(\rbzero.spi_registers.spi_cmd[2] ),
    .Y(_02581_));
 sky130_fd_sc_hd__and4b_1 _18867_ (.A_N(\rbzero.spi_registers.spi_cmd[3] ),
    .B(_02581_),
    .C(\rbzero.spi_registers.spi_cmd[1] ),
    .D(\rbzero.spi_registers.spi_cmd[0] ),
    .X(_02582_));
 sky130_fd_sc_hd__xnor2_1 _18868_ (.A(\rbzero.spi_registers.spi_counter[1] ),
    .B(_02582_),
    .Y(_02583_));
 sky130_fd_sc_hd__o21a_1 _18869_ (.A1(\rbzero.spi_registers.spi_counter[3] ),
    .A2(_02579_),
    .B1(_02583_),
    .X(_02584_));
 sky130_fd_sc_hd__a21o_1 _18870_ (.A1(\rbzero.spi_registers.spi_cmd[1] ),
    .A2(\rbzero.spi_registers.spi_cmd[0] ),
    .B1(_02579_),
    .X(_02585_));
 sky130_fd_sc_hd__xnor2_1 _18871_ (.A(\rbzero.spi_registers.spi_counter[2] ),
    .B(_02585_),
    .Y(_02586_));
 sky130_fd_sc_hd__and4bb_1 _18872_ (.A_N(_02577_),
    .B_N(_02580_),
    .C(_02584_),
    .D(_02586_),
    .X(_02587_));
 sky130_fd_sc_hd__o21ai_1 _18873_ (.A1(\rbzero.spi_registers.spi_counter[0] ),
    .A2(_02587_),
    .B1(_02576_),
    .Y(_02588_));
 sky130_fd_sc_hd__nor2_2 _18874_ (.A(\rbzero.spi_registers.ss_buffer[1] ),
    .B(_03442_),
    .Y(_02589_));
 sky130_fd_sc_hd__o211a_1 _18875_ (.A1(\rbzero.spi_registers.spi_counter[0] ),
    .A2(_02576_),
    .B1(_02588_),
    .C1(_02589_),
    .X(_00629_));
 sky130_fd_sc_hd__a21boi_1 _18876_ (.A1(_02576_),
    .A2(_02587_),
    .B1_N(_02589_),
    .Y(_02590_));
 sky130_fd_sc_hd__nand3_1 _18877_ (.A(\rbzero.spi_registers.spi_counter[1] ),
    .B(\rbzero.spi_registers.spi_counter[0] ),
    .C(_02576_),
    .Y(_02591_));
 sky130_fd_sc_hd__a21o_1 _18878_ (.A1(\rbzero.spi_registers.spi_counter[0] ),
    .A2(_02576_),
    .B1(\rbzero.spi_registers.spi_counter[1] ),
    .X(_02592_));
 sky130_fd_sc_hd__and3_1 _18879_ (.A(_02590_),
    .B(_02591_),
    .C(_02592_),
    .X(_02593_));
 sky130_fd_sc_hd__clkbuf_1 _18880_ (.A(_02593_),
    .X(_00630_));
 sky130_fd_sc_hd__and4_1 _18881_ (.A(\rbzero.spi_registers.spi_counter[2] ),
    .B(\rbzero.spi_registers.spi_counter[1] ),
    .C(\rbzero.spi_registers.spi_counter[0] ),
    .D(_02576_),
    .X(_02594_));
 sky130_fd_sc_hd__a31o_1 _18882_ (.A1(\rbzero.spi_registers.spi_counter[1] ),
    .A2(\rbzero.spi_registers.spi_counter[0] ),
    .A3(_02576_),
    .B1(\rbzero.spi_registers.spi_counter[2] ),
    .X(_02595_));
 sky130_fd_sc_hd__and3b_1 _18883_ (.A_N(_02594_),
    .B(_02595_),
    .C(_02590_),
    .X(_02596_));
 sky130_fd_sc_hd__clkbuf_1 _18884_ (.A(_02596_),
    .X(_00631_));
 sky130_fd_sc_hd__nand2_1 _18885_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(_02594_),
    .Y(_02597_));
 sky130_fd_sc_hd__or2_1 _18886_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(_02594_),
    .X(_02598_));
 sky130_fd_sc_hd__and3_1 _18887_ (.A(_02590_),
    .B(_02597_),
    .C(_02598_),
    .X(_02599_));
 sky130_fd_sc_hd__clkbuf_1 _18888_ (.A(_02599_),
    .X(_00632_));
 sky130_fd_sc_hd__xnor2_1 _18889_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(_02597_),
    .Y(_02600_));
 sky130_fd_sc_hd__and2_1 _18890_ (.A(_02590_),
    .B(_02600_),
    .X(_02601_));
 sky130_fd_sc_hd__clkbuf_1 _18891_ (.A(_02601_),
    .X(_00633_));
 sky130_fd_sc_hd__and4_1 _18892_ (.A(\rbzero.spi_registers.spi_counter[5] ),
    .B(\rbzero.spi_registers.spi_counter[4] ),
    .C(\rbzero.spi_registers.spi_counter[3] ),
    .D(_02594_),
    .X(_02602_));
 sky130_fd_sc_hd__a31o_1 _18893_ (.A1(\rbzero.spi_registers.spi_counter[4] ),
    .A2(\rbzero.spi_registers.spi_counter[3] ),
    .A3(_02594_),
    .B1(\rbzero.spi_registers.spi_counter[5] ),
    .X(_02603_));
 sky130_fd_sc_hd__and3b_1 _18894_ (.A_N(_02602_),
    .B(_02589_),
    .C(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__clkbuf_1 _18895_ (.A(_02604_),
    .X(_00634_));
 sky130_fd_sc_hd__o21ai_1 _18896_ (.A1(\rbzero.spi_registers.spi_counter[6] ),
    .A2(_02602_),
    .B1(_02589_),
    .Y(_02605_));
 sky130_fd_sc_hd__a21oi_1 _18897_ (.A1(\rbzero.spi_registers.spi_counter[6] ),
    .A2(_02602_),
    .B1(_02605_),
    .Y(_00635_));
 sky130_fd_sc_hd__nand2_2 _18898_ (.A(\rbzero.pov.spi_done ),
    .B(_03292_),
    .Y(_02606_));
 sky130_fd_sc_hd__clkbuf_4 _18899_ (.A(_02606_),
    .X(_02607_));
 sky130_fd_sc_hd__clkbuf_4 _18900_ (.A(_02607_),
    .X(_02608_));
 sky130_fd_sc_hd__mux2_1 _18901_ (.A0(\rbzero.pov.spi_buffer[0] ),
    .A1(\rbzero.pov.ready_buffer[0] ),
    .S(_02608_),
    .X(_02609_));
 sky130_fd_sc_hd__clkbuf_1 _18902_ (.A(_02609_),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _18903_ (.A0(\rbzero.pov.spi_buffer[1] ),
    .A1(\rbzero.pov.ready_buffer[1] ),
    .S(_02608_),
    .X(_02610_));
 sky130_fd_sc_hd__clkbuf_1 _18904_ (.A(_02610_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _18905_ (.A0(\rbzero.pov.spi_buffer[2] ),
    .A1(\rbzero.pov.ready_buffer[2] ),
    .S(_02608_),
    .X(_02611_));
 sky130_fd_sc_hd__clkbuf_1 _18906_ (.A(_02611_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _18907_ (.A0(\rbzero.pov.spi_buffer[3] ),
    .A1(\rbzero.pov.ready_buffer[3] ),
    .S(_02608_),
    .X(_02612_));
 sky130_fd_sc_hd__clkbuf_1 _18908_ (.A(_02612_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _18909_ (.A0(\rbzero.pov.spi_buffer[4] ),
    .A1(\rbzero.pov.ready_buffer[4] ),
    .S(_02608_),
    .X(_02613_));
 sky130_fd_sc_hd__clkbuf_1 _18910_ (.A(_02613_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _18911_ (.A0(\rbzero.pov.spi_buffer[5] ),
    .A1(\rbzero.pov.ready_buffer[5] ),
    .S(_02608_),
    .X(_02614_));
 sky130_fd_sc_hd__clkbuf_1 _18912_ (.A(_02614_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _18913_ (.A0(\rbzero.pov.spi_buffer[6] ),
    .A1(\rbzero.pov.ready_buffer[6] ),
    .S(_02608_),
    .X(_02615_));
 sky130_fd_sc_hd__clkbuf_1 _18914_ (.A(_02615_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _18915_ (.A0(\rbzero.pov.spi_buffer[7] ),
    .A1(\rbzero.pov.ready_buffer[7] ),
    .S(_02608_),
    .X(_02616_));
 sky130_fd_sc_hd__clkbuf_1 _18916_ (.A(_02616_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _18917_ (.A0(\rbzero.pov.spi_buffer[8] ),
    .A1(\rbzero.pov.ready_buffer[8] ),
    .S(_02608_),
    .X(_02617_));
 sky130_fd_sc_hd__clkbuf_1 _18918_ (.A(_02617_),
    .X(_00644_));
 sky130_fd_sc_hd__clkbuf_4 _18919_ (.A(_02607_),
    .X(_02618_));
 sky130_fd_sc_hd__mux2_1 _18920_ (.A0(\rbzero.pov.spi_buffer[9] ),
    .A1(\rbzero.pov.ready_buffer[9] ),
    .S(_02618_),
    .X(_02619_));
 sky130_fd_sc_hd__clkbuf_1 _18921_ (.A(_02619_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _18922_ (.A0(\rbzero.pov.spi_buffer[10] ),
    .A1(\rbzero.pov.ready_buffer[10] ),
    .S(_02618_),
    .X(_02620_));
 sky130_fd_sc_hd__clkbuf_1 _18923_ (.A(_02620_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _18924_ (.A0(\rbzero.pov.spi_buffer[11] ),
    .A1(\rbzero.pov.ready_buffer[11] ),
    .S(_02618_),
    .X(_02621_));
 sky130_fd_sc_hd__clkbuf_1 _18925_ (.A(_02621_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _18926_ (.A0(\rbzero.pov.spi_buffer[12] ),
    .A1(\rbzero.pov.ready_buffer[12] ),
    .S(_02618_),
    .X(_02622_));
 sky130_fd_sc_hd__clkbuf_1 _18927_ (.A(_02622_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _18928_ (.A0(\rbzero.pov.spi_buffer[13] ),
    .A1(\rbzero.pov.ready_buffer[13] ),
    .S(_02618_),
    .X(_02623_));
 sky130_fd_sc_hd__clkbuf_1 _18929_ (.A(_02623_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _18930_ (.A0(\rbzero.pov.spi_buffer[14] ),
    .A1(\rbzero.pov.ready_buffer[14] ),
    .S(_02618_),
    .X(_02624_));
 sky130_fd_sc_hd__clkbuf_1 _18931_ (.A(_02624_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _18932_ (.A0(\rbzero.pov.spi_buffer[15] ),
    .A1(\rbzero.pov.ready_buffer[15] ),
    .S(_02618_),
    .X(_02625_));
 sky130_fd_sc_hd__clkbuf_1 _18933_ (.A(_02625_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _18934_ (.A0(\rbzero.pov.spi_buffer[16] ),
    .A1(\rbzero.pov.ready_buffer[16] ),
    .S(_02618_),
    .X(_02626_));
 sky130_fd_sc_hd__clkbuf_1 _18935_ (.A(_02626_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _18936_ (.A0(\rbzero.pov.spi_buffer[17] ),
    .A1(\rbzero.pov.ready_buffer[17] ),
    .S(_02618_),
    .X(_02627_));
 sky130_fd_sc_hd__clkbuf_1 _18937_ (.A(_02627_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _18938_ (.A0(\rbzero.pov.spi_buffer[18] ),
    .A1(\rbzero.pov.ready_buffer[18] ),
    .S(_02618_),
    .X(_02628_));
 sky130_fd_sc_hd__clkbuf_1 _18939_ (.A(_02628_),
    .X(_00654_));
 sky130_fd_sc_hd__clkbuf_4 _18940_ (.A(_02607_),
    .X(_02629_));
 sky130_fd_sc_hd__mux2_1 _18941_ (.A0(\rbzero.pov.spi_buffer[19] ),
    .A1(\rbzero.pov.ready_buffer[19] ),
    .S(_02629_),
    .X(_02630_));
 sky130_fd_sc_hd__clkbuf_1 _18942_ (.A(_02630_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _18943_ (.A0(\rbzero.pov.spi_buffer[20] ),
    .A1(\rbzero.pov.ready_buffer[20] ),
    .S(_02629_),
    .X(_02631_));
 sky130_fd_sc_hd__clkbuf_1 _18944_ (.A(_02631_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _18945_ (.A0(\rbzero.pov.spi_buffer[21] ),
    .A1(\rbzero.pov.ready_buffer[21] ),
    .S(_02629_),
    .X(_02632_));
 sky130_fd_sc_hd__clkbuf_1 _18946_ (.A(_02632_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _18947_ (.A0(\rbzero.pov.spi_buffer[22] ),
    .A1(\rbzero.pov.ready_buffer[22] ),
    .S(_02629_),
    .X(_02633_));
 sky130_fd_sc_hd__clkbuf_1 _18948_ (.A(_02633_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _18949_ (.A0(\rbzero.pov.spi_buffer[23] ),
    .A1(\rbzero.pov.ready_buffer[23] ),
    .S(_02629_),
    .X(_02634_));
 sky130_fd_sc_hd__clkbuf_1 _18950_ (.A(_02634_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _18951_ (.A0(\rbzero.pov.spi_buffer[24] ),
    .A1(\rbzero.pov.ready_buffer[24] ),
    .S(_02629_),
    .X(_02635_));
 sky130_fd_sc_hd__clkbuf_1 _18952_ (.A(_02635_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _18953_ (.A0(\rbzero.pov.spi_buffer[25] ),
    .A1(\rbzero.pov.ready_buffer[25] ),
    .S(_02629_),
    .X(_02636_));
 sky130_fd_sc_hd__clkbuf_1 _18954_ (.A(_02636_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _18955_ (.A0(\rbzero.pov.spi_buffer[26] ),
    .A1(\rbzero.pov.ready_buffer[26] ),
    .S(_02629_),
    .X(_02637_));
 sky130_fd_sc_hd__clkbuf_1 _18956_ (.A(_02637_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _18957_ (.A0(\rbzero.pov.spi_buffer[27] ),
    .A1(\rbzero.pov.ready_buffer[27] ),
    .S(_02629_),
    .X(_02638_));
 sky130_fd_sc_hd__clkbuf_1 _18958_ (.A(_02638_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _18959_ (.A0(\rbzero.pov.spi_buffer[28] ),
    .A1(\rbzero.pov.ready_buffer[28] ),
    .S(_02629_),
    .X(_02639_));
 sky130_fd_sc_hd__clkbuf_1 _18960_ (.A(_02639_),
    .X(_00664_));
 sky130_fd_sc_hd__clkbuf_4 _18961_ (.A(_02607_),
    .X(_02640_));
 sky130_fd_sc_hd__mux2_1 _18962_ (.A0(\rbzero.pov.spi_buffer[29] ),
    .A1(\rbzero.pov.ready_buffer[29] ),
    .S(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__clkbuf_1 _18963_ (.A(_02641_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _18964_ (.A0(\rbzero.pov.spi_buffer[30] ),
    .A1(\rbzero.pov.ready_buffer[30] ),
    .S(_02640_),
    .X(_02642_));
 sky130_fd_sc_hd__clkbuf_1 _18965_ (.A(_02642_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _18966_ (.A0(\rbzero.pov.spi_buffer[31] ),
    .A1(\rbzero.pov.ready_buffer[31] ),
    .S(_02640_),
    .X(_02643_));
 sky130_fd_sc_hd__clkbuf_1 _18967_ (.A(_02643_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _18968_ (.A0(\rbzero.pov.spi_buffer[32] ),
    .A1(\rbzero.pov.ready_buffer[32] ),
    .S(_02640_),
    .X(_02644_));
 sky130_fd_sc_hd__clkbuf_1 _18969_ (.A(_02644_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _18970_ (.A0(\rbzero.pov.spi_buffer[33] ),
    .A1(\rbzero.pov.ready_buffer[33] ),
    .S(_02640_),
    .X(_02645_));
 sky130_fd_sc_hd__clkbuf_1 _18971_ (.A(_02645_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _18972_ (.A0(\rbzero.pov.spi_buffer[34] ),
    .A1(\rbzero.pov.ready_buffer[34] ),
    .S(_02640_),
    .X(_02646_));
 sky130_fd_sc_hd__clkbuf_1 _18973_ (.A(_02646_),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _18974_ (.A0(\rbzero.pov.spi_buffer[35] ),
    .A1(\rbzero.pov.ready_buffer[35] ),
    .S(_02640_),
    .X(_02647_));
 sky130_fd_sc_hd__clkbuf_1 _18975_ (.A(_02647_),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _18976_ (.A0(\rbzero.pov.spi_buffer[36] ),
    .A1(\rbzero.pov.ready_buffer[36] ),
    .S(_02640_),
    .X(_02648_));
 sky130_fd_sc_hd__clkbuf_1 _18977_ (.A(_02648_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _18978_ (.A0(\rbzero.pov.spi_buffer[37] ),
    .A1(\rbzero.pov.ready_buffer[37] ),
    .S(_02640_),
    .X(_02649_));
 sky130_fd_sc_hd__clkbuf_1 _18979_ (.A(_02649_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _18980_ (.A0(\rbzero.pov.spi_buffer[38] ),
    .A1(\rbzero.pov.ready_buffer[38] ),
    .S(_02640_),
    .X(_02650_));
 sky130_fd_sc_hd__clkbuf_1 _18981_ (.A(_02650_),
    .X(_00674_));
 sky130_fd_sc_hd__clkbuf_4 _18982_ (.A(_02607_),
    .X(_02651_));
 sky130_fd_sc_hd__mux2_1 _18983_ (.A0(\rbzero.pov.spi_buffer[39] ),
    .A1(\rbzero.pov.ready_buffer[39] ),
    .S(_02651_),
    .X(_02652_));
 sky130_fd_sc_hd__clkbuf_1 _18984_ (.A(_02652_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _18985_ (.A0(\rbzero.pov.spi_buffer[40] ),
    .A1(\rbzero.pov.ready_buffer[40] ),
    .S(_02651_),
    .X(_02653_));
 sky130_fd_sc_hd__clkbuf_1 _18986_ (.A(_02653_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _18987_ (.A0(\rbzero.pov.spi_buffer[41] ),
    .A1(\rbzero.pov.ready_buffer[41] ),
    .S(_02651_),
    .X(_02654_));
 sky130_fd_sc_hd__clkbuf_1 _18988_ (.A(_02654_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _18989_ (.A0(\rbzero.pov.spi_buffer[42] ),
    .A1(\rbzero.pov.ready_buffer[42] ),
    .S(_02651_),
    .X(_02655_));
 sky130_fd_sc_hd__clkbuf_1 _18990_ (.A(_02655_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _18991_ (.A0(\rbzero.pov.spi_buffer[43] ),
    .A1(\rbzero.pov.ready_buffer[43] ),
    .S(_02651_),
    .X(_02656_));
 sky130_fd_sc_hd__clkbuf_1 _18992_ (.A(_02656_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _18993_ (.A0(\rbzero.pov.spi_buffer[44] ),
    .A1(\rbzero.pov.ready_buffer[44] ),
    .S(_02651_),
    .X(_02657_));
 sky130_fd_sc_hd__clkbuf_1 _18994_ (.A(_02657_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _18995_ (.A0(\rbzero.pov.spi_buffer[45] ),
    .A1(\rbzero.pov.ready_buffer[45] ),
    .S(_02651_),
    .X(_02658_));
 sky130_fd_sc_hd__clkbuf_1 _18996_ (.A(_02658_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _18997_ (.A0(\rbzero.pov.spi_buffer[46] ),
    .A1(\rbzero.pov.ready_buffer[46] ),
    .S(_02651_),
    .X(_02659_));
 sky130_fd_sc_hd__clkbuf_1 _18998_ (.A(_02659_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _18999_ (.A0(\rbzero.pov.spi_buffer[47] ),
    .A1(\rbzero.pov.ready_buffer[47] ),
    .S(_02651_),
    .X(_02660_));
 sky130_fd_sc_hd__clkbuf_1 _19000_ (.A(_02660_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _19001_ (.A0(\rbzero.pov.spi_buffer[48] ),
    .A1(\rbzero.pov.ready_buffer[48] ),
    .S(_02651_),
    .X(_02661_));
 sky130_fd_sc_hd__clkbuf_1 _19002_ (.A(_02661_),
    .X(_00684_));
 sky130_fd_sc_hd__clkbuf_4 _19003_ (.A(_02606_),
    .X(_02662_));
 sky130_fd_sc_hd__mux2_1 _19004_ (.A0(\rbzero.pov.spi_buffer[49] ),
    .A1(\rbzero.pov.ready_buffer[49] ),
    .S(_02662_),
    .X(_02663_));
 sky130_fd_sc_hd__clkbuf_1 _19005_ (.A(_02663_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _19006_ (.A0(\rbzero.pov.spi_buffer[50] ),
    .A1(\rbzero.pov.ready_buffer[50] ),
    .S(_02662_),
    .X(_02664_));
 sky130_fd_sc_hd__clkbuf_1 _19007_ (.A(_02664_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _19008_ (.A0(\rbzero.pov.spi_buffer[51] ),
    .A1(\rbzero.pov.ready_buffer[51] ),
    .S(_02662_),
    .X(_02665_));
 sky130_fd_sc_hd__clkbuf_1 _19009_ (.A(_02665_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _19010_ (.A0(\rbzero.pov.spi_buffer[52] ),
    .A1(\rbzero.pov.ready_buffer[52] ),
    .S(_02662_),
    .X(_02666_));
 sky130_fd_sc_hd__clkbuf_1 _19011_ (.A(_02666_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _19012_ (.A0(\rbzero.pov.spi_buffer[53] ),
    .A1(\rbzero.pov.ready_buffer[53] ),
    .S(_02662_),
    .X(_02667_));
 sky130_fd_sc_hd__clkbuf_1 _19013_ (.A(_02667_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _19014_ (.A0(\rbzero.pov.spi_buffer[54] ),
    .A1(\rbzero.pov.ready_buffer[54] ),
    .S(_02662_),
    .X(_02668_));
 sky130_fd_sc_hd__clkbuf_1 _19015_ (.A(_02668_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _19016_ (.A0(\rbzero.pov.spi_buffer[55] ),
    .A1(\rbzero.pov.ready_buffer[55] ),
    .S(_02662_),
    .X(_02669_));
 sky130_fd_sc_hd__clkbuf_1 _19017_ (.A(_02669_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _19018_ (.A0(\rbzero.pov.spi_buffer[56] ),
    .A1(\rbzero.pov.ready_buffer[56] ),
    .S(_02662_),
    .X(_02670_));
 sky130_fd_sc_hd__clkbuf_1 _19019_ (.A(_02670_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _19020_ (.A0(\rbzero.pov.spi_buffer[57] ),
    .A1(\rbzero.pov.ready_buffer[57] ),
    .S(_02662_),
    .X(_02671_));
 sky130_fd_sc_hd__clkbuf_1 _19021_ (.A(_02671_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _19022_ (.A0(\rbzero.pov.spi_buffer[58] ),
    .A1(\rbzero.pov.ready_buffer[58] ),
    .S(_02662_),
    .X(_02672_));
 sky130_fd_sc_hd__clkbuf_1 _19023_ (.A(_02672_),
    .X(_00694_));
 sky130_fd_sc_hd__clkbuf_4 _19024_ (.A(_02606_),
    .X(_02673_));
 sky130_fd_sc_hd__mux2_1 _19025_ (.A0(\rbzero.pov.spi_buffer[59] ),
    .A1(\rbzero.pov.ready_buffer[59] ),
    .S(_02673_),
    .X(_02674_));
 sky130_fd_sc_hd__clkbuf_1 _19026_ (.A(_02674_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _19027_ (.A0(\rbzero.pov.spi_buffer[60] ),
    .A1(\rbzero.pov.ready_buffer[60] ),
    .S(_02673_),
    .X(_02675_));
 sky130_fd_sc_hd__clkbuf_1 _19028_ (.A(_02675_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _19029_ (.A0(\rbzero.pov.spi_buffer[61] ),
    .A1(\rbzero.pov.ready_buffer[61] ),
    .S(_02673_),
    .X(_02676_));
 sky130_fd_sc_hd__clkbuf_1 _19030_ (.A(_02676_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _19031_ (.A0(\rbzero.pov.spi_buffer[62] ),
    .A1(\rbzero.pov.ready_buffer[62] ),
    .S(_02673_),
    .X(_02677_));
 sky130_fd_sc_hd__clkbuf_1 _19032_ (.A(_02677_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _19033_ (.A0(\rbzero.pov.spi_buffer[63] ),
    .A1(\rbzero.pov.ready_buffer[63] ),
    .S(_02673_),
    .X(_02678_));
 sky130_fd_sc_hd__clkbuf_1 _19034_ (.A(_02678_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _19035_ (.A0(\rbzero.pov.spi_buffer[64] ),
    .A1(\rbzero.pov.ready_buffer[64] ),
    .S(_02673_),
    .X(_02679_));
 sky130_fd_sc_hd__clkbuf_1 _19036_ (.A(_02679_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _19037_ (.A0(\rbzero.pov.spi_buffer[65] ),
    .A1(\rbzero.pov.ready_buffer[65] ),
    .S(_02673_),
    .X(_02680_));
 sky130_fd_sc_hd__clkbuf_1 _19038_ (.A(_02680_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _19039_ (.A0(\rbzero.pov.spi_buffer[66] ),
    .A1(\rbzero.pov.ready_buffer[66] ),
    .S(_02673_),
    .X(_02681_));
 sky130_fd_sc_hd__clkbuf_1 _19040_ (.A(_02681_),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _19041_ (.A0(\rbzero.pov.spi_buffer[67] ),
    .A1(\rbzero.pov.ready_buffer[67] ),
    .S(_02673_),
    .X(_02682_));
 sky130_fd_sc_hd__clkbuf_1 _19042_ (.A(_02682_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _19043_ (.A0(\rbzero.pov.spi_buffer[68] ),
    .A1(\rbzero.pov.ready_buffer[68] ),
    .S(_02673_),
    .X(_02683_));
 sky130_fd_sc_hd__clkbuf_1 _19044_ (.A(_02683_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _19045_ (.A0(\rbzero.pov.spi_buffer[69] ),
    .A1(\rbzero.pov.ready_buffer[69] ),
    .S(_02607_),
    .X(_02684_));
 sky130_fd_sc_hd__clkbuf_1 _19046_ (.A(_02684_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _19047_ (.A0(\rbzero.pov.spi_buffer[70] ),
    .A1(\rbzero.pov.ready_buffer[70] ),
    .S(_02607_),
    .X(_02685_));
 sky130_fd_sc_hd__clkbuf_1 _19048_ (.A(_02685_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _19049_ (.A0(\rbzero.pov.spi_buffer[71] ),
    .A1(\rbzero.pov.ready_buffer[71] ),
    .S(_02607_),
    .X(_02686_));
 sky130_fd_sc_hd__clkbuf_1 _19050_ (.A(_02686_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _19051_ (.A0(\rbzero.pov.spi_buffer[72] ),
    .A1(\rbzero.pov.ready_buffer[72] ),
    .S(_02607_),
    .X(_02687_));
 sky130_fd_sc_hd__clkbuf_1 _19052_ (.A(_02687_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _19053_ (.A0(\rbzero.pov.spi_buffer[73] ),
    .A1(\rbzero.pov.ready_buffer[73] ),
    .S(_02607_),
    .X(_02688_));
 sky130_fd_sc_hd__clkbuf_1 _19054_ (.A(_02688_),
    .X(_00709_));
 sky130_fd_sc_hd__o311a_1 _19055_ (.A1(\rbzero.spi_registers.spi_counter[3] ),
    .A2(\rbzero.spi_registers.spi_counter[2] ),
    .A3(_02577_),
    .B1(_02576_),
    .C1(_02589_),
    .X(_02689_));
 sky130_fd_sc_hd__clkbuf_4 _19056_ (.A(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__mux2_1 _19057_ (.A0(\rbzero.spi_registers.spi_buffer[0] ),
    .A1(\rbzero.spi_registers.mosi ),
    .S(_02690_),
    .X(_02691_));
 sky130_fd_sc_hd__clkbuf_1 _19058_ (.A(_02691_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _19059_ (.A0(\rbzero.spi_registers.spi_buffer[1] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_02690_),
    .X(_02692_));
 sky130_fd_sc_hd__clkbuf_1 _19060_ (.A(_02692_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _19061_ (.A0(\rbzero.spi_registers.spi_buffer[2] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_02690_),
    .X(_02693_));
 sky130_fd_sc_hd__clkbuf_1 _19062_ (.A(_02693_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _19063_ (.A0(\rbzero.spi_registers.spi_buffer[3] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_02690_),
    .X(_02694_));
 sky130_fd_sc_hd__clkbuf_1 _19064_ (.A(_02694_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _19065_ (.A0(\rbzero.spi_registers.spi_buffer[4] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_02690_),
    .X(_02695_));
 sky130_fd_sc_hd__clkbuf_1 _19066_ (.A(_02695_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _19067_ (.A0(\rbzero.spi_registers.spi_buffer[5] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_02690_),
    .X(_02696_));
 sky130_fd_sc_hd__clkbuf_1 _19068_ (.A(_02696_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _19069_ (.A0(\rbzero.spi_registers.spi_buffer[6] ),
    .A1(\rbzero.spi_registers.spi_buffer[5] ),
    .S(_02690_),
    .X(_02697_));
 sky130_fd_sc_hd__clkbuf_1 _19070_ (.A(_02697_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _19071_ (.A0(\rbzero.spi_registers.spi_buffer[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_02690_),
    .X(_02698_));
 sky130_fd_sc_hd__clkbuf_1 _19072_ (.A(_02698_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _19073_ (.A0(\rbzero.spi_registers.spi_buffer[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_02690_),
    .X(_02699_));
 sky130_fd_sc_hd__clkbuf_1 _19074_ (.A(_02699_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _19075_ (.A0(\rbzero.spi_registers.spi_buffer[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_02690_),
    .X(_02700_));
 sky130_fd_sc_hd__clkbuf_1 _19076_ (.A(_02700_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _19077_ (.A0(\rbzero.spi_registers.spi_buffer[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_02689_),
    .X(_02701_));
 sky130_fd_sc_hd__clkbuf_1 _19078_ (.A(_02701_),
    .X(_00720_));
 sky130_fd_sc_hd__nand2_1 _19079_ (.A(_02589_),
    .B(_02576_),
    .Y(_02702_));
 sky130_fd_sc_hd__or4_2 _19080_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(\rbzero.spi_registers.spi_counter[2] ),
    .C(_02577_),
    .D(_02702_),
    .X(_02703_));
 sky130_fd_sc_hd__mux2_1 _19081_ (.A0(\rbzero.spi_registers.mosi ),
    .A1(\rbzero.spi_registers.spi_cmd[0] ),
    .S(_02703_),
    .X(_02704_));
 sky130_fd_sc_hd__clkbuf_1 _19082_ (.A(_02704_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _19083_ (.A0(\rbzero.spi_registers.spi_cmd[0] ),
    .A1(\rbzero.spi_registers.spi_cmd[1] ),
    .S(_02703_),
    .X(_02705_));
 sky130_fd_sc_hd__clkbuf_1 _19084_ (.A(_02705_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _19085_ (.A0(\rbzero.spi_registers.spi_cmd[1] ),
    .A1(\rbzero.spi_registers.spi_cmd[2] ),
    .S(_02703_),
    .X(_02706_));
 sky130_fd_sc_hd__clkbuf_1 _19086_ (.A(_02706_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _19087_ (.A0(\rbzero.spi_registers.spi_cmd[2] ),
    .A1(\rbzero.spi_registers.spi_cmd[3] ),
    .S(_02703_),
    .X(_02707_));
 sky130_fd_sc_hd__clkbuf_1 _19088_ (.A(_02707_),
    .X(_00724_));
 sky130_fd_sc_hd__buf_6 _19089_ (.A(_03442_),
    .X(_02708_));
 sky130_fd_sc_hd__mux2_1 _19090_ (.A0(net43),
    .A1(\rbzero.spi_registers.mosi_buffer[0] ),
    .S(_02708_),
    .X(_02709_));
 sky130_fd_sc_hd__clkbuf_1 _19091_ (.A(_02709_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _19092_ (.A0(\rbzero.spi_registers.mosi ),
    .A1(\rbzero.spi_registers.mosi_buffer[0] ),
    .S(_04920_),
    .X(_02710_));
 sky130_fd_sc_hd__clkbuf_1 _19093_ (.A(_02710_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _19094_ (.A0(net42),
    .A1(\rbzero.spi_registers.ss_buffer[0] ),
    .S(_02708_),
    .X(_02711_));
 sky130_fd_sc_hd__clkbuf_1 _19095_ (.A(_02711_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _19096_ (.A0(\rbzero.spi_registers.ss_buffer[1] ),
    .A1(\rbzero.spi_registers.ss_buffer[0] ),
    .S(_04920_),
    .X(_02712_));
 sky130_fd_sc_hd__clkbuf_1 _19097_ (.A(_02712_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _19098_ (.A0(net44),
    .A1(\rbzero.spi_registers.sclk_buffer[0] ),
    .S(_02708_),
    .X(_02713_));
 sky130_fd_sc_hd__clkbuf_1 _19099_ (.A(_02713_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _19100_ (.A0(\rbzero.spi_registers.sclk_buffer[1] ),
    .A1(\rbzero.spi_registers.sclk_buffer[0] ),
    .S(_09243_),
    .X(_02714_));
 sky130_fd_sc_hd__clkbuf_1 _19101_ (.A(_02714_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _19102_ (.A0(\rbzero.spi_registers.sclk_buffer[2] ),
    .A1(\rbzero.spi_registers.sclk_buffer[1] ),
    .S(_09243_),
    .X(_02715_));
 sky130_fd_sc_hd__clkbuf_1 _19103_ (.A(_02715_),
    .X(_00731_));
 sky130_fd_sc_hd__and3_1 _19104_ (.A(\gpout0.vpos[2] ),
    .B(\gpout0.vpos[1] ),
    .C(\gpout0.vpos[0] ),
    .X(_02716_));
 sky130_fd_sc_hd__inv_2 _19105_ (.A(_02716_),
    .Y(_02717_));
 sky130_fd_sc_hd__nor2_1 _19106_ (.A(_04246_),
    .B(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__and2_1 _19107_ (.A(_03808_),
    .B(_02718_),
    .X(_02719_));
 sky130_fd_sc_hd__and4_4 _19108_ (.A(_04111_),
    .B(_04252_),
    .C(_04113_),
    .D(_02719_),
    .X(_02720_));
 sky130_fd_sc_hd__buf_4 _19109_ (.A(_02720_),
    .X(_02721_));
 sky130_fd_sc_hd__and2_1 _19110_ (.A(\rbzero.spi_registers.got_new_other ),
    .B(_02721_),
    .X(_02722_));
 sky130_fd_sc_hd__buf_2 _19111_ (.A(_02722_),
    .X(_02723_));
 sky130_fd_sc_hd__clkbuf_4 _19112_ (.A(_02721_),
    .X(_02724_));
 sky130_fd_sc_hd__nand2_2 _19113_ (.A(\rbzero.spi_registers.got_new_other ),
    .B(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__or2_1 _19114_ (.A(\rbzero.spi_registers.new_other[6] ),
    .B(_02725_),
    .X(_02726_));
 sky130_fd_sc_hd__buf_4 _19115_ (.A(_09243_),
    .X(_02727_));
 sky130_fd_sc_hd__clkbuf_4 _19116_ (.A(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__o211a_1 _19117_ (.A1(\rbzero.otherx[0] ),
    .A2(_02723_),
    .B1(_02726_),
    .C1(_02728_),
    .X(_00732_));
 sky130_fd_sc_hd__or2_1 _19118_ (.A(\rbzero.spi_registers.new_other[7] ),
    .B(_02725_),
    .X(_02729_));
 sky130_fd_sc_hd__o211a_1 _19119_ (.A1(\rbzero.otherx[1] ),
    .A2(_02723_),
    .B1(_02729_),
    .C1(_02728_),
    .X(_00733_));
 sky130_fd_sc_hd__or2_1 _19120_ (.A(\rbzero.spi_registers.new_other[8] ),
    .B(_02725_),
    .X(_02730_));
 sky130_fd_sc_hd__o211a_1 _19121_ (.A1(\rbzero.otherx[2] ),
    .A2(_02723_),
    .B1(_02730_),
    .C1(_02728_),
    .X(_00734_));
 sky130_fd_sc_hd__or2_1 _19122_ (.A(\rbzero.spi_registers.new_other[9] ),
    .B(_02725_),
    .X(_02731_));
 sky130_fd_sc_hd__o211a_1 _19123_ (.A1(\rbzero.otherx[3] ),
    .A2(_02723_),
    .B1(_02731_),
    .C1(_02728_),
    .X(_00735_));
 sky130_fd_sc_hd__or2_1 _19124_ (.A(\rbzero.spi_registers.new_other[10] ),
    .B(_02725_),
    .X(_02732_));
 sky130_fd_sc_hd__o211a_1 _19125_ (.A1(\rbzero.otherx[4] ),
    .A2(_02723_),
    .B1(_02732_),
    .C1(_02728_),
    .X(_00736_));
 sky130_fd_sc_hd__or2_1 _19126_ (.A(\rbzero.spi_registers.new_other[0] ),
    .B(_02725_),
    .X(_02733_));
 sky130_fd_sc_hd__o211a_1 _19127_ (.A1(\rbzero.othery[0] ),
    .A2(_02723_),
    .B1(_02733_),
    .C1(_02728_),
    .X(_00737_));
 sky130_fd_sc_hd__or2_1 _19128_ (.A(\rbzero.spi_registers.new_other[1] ),
    .B(_02725_),
    .X(_02734_));
 sky130_fd_sc_hd__o211a_1 _19129_ (.A1(\rbzero.othery[1] ),
    .A2(_02723_),
    .B1(_02734_),
    .C1(_02728_),
    .X(_00738_));
 sky130_fd_sc_hd__or2_1 _19130_ (.A(\rbzero.spi_registers.new_other[2] ),
    .B(_02725_),
    .X(_02735_));
 sky130_fd_sc_hd__o211a_1 _19131_ (.A1(\rbzero.othery[2] ),
    .A2(_02723_),
    .B1(_02735_),
    .C1(_02728_),
    .X(_00739_));
 sky130_fd_sc_hd__or2_1 _19132_ (.A(\rbzero.spi_registers.new_other[3] ),
    .B(_02725_),
    .X(_02736_));
 sky130_fd_sc_hd__o211a_1 _19133_ (.A1(\rbzero.othery[3] ),
    .A2(_02723_),
    .B1(_02736_),
    .C1(_02728_),
    .X(_00740_));
 sky130_fd_sc_hd__or2_1 _19134_ (.A(\rbzero.spi_registers.new_other[4] ),
    .B(_02725_),
    .X(_02737_));
 sky130_fd_sc_hd__buf_2 _19135_ (.A(_02727_),
    .X(_02738_));
 sky130_fd_sc_hd__o211a_1 _19136_ (.A1(\rbzero.othery[4] ),
    .A2(_02723_),
    .B1(_02737_),
    .C1(_02738_),
    .X(_00741_));
 sky130_fd_sc_hd__inv_2 _19137_ (.A(\rbzero.spi_registers.got_new_vinf ),
    .Y(_02739_));
 sky130_fd_sc_hd__nand4_4 _19138_ (.A(_04111_),
    .B(_04252_),
    .C(_04113_),
    .D(_02719_),
    .Y(_02740_));
 sky130_fd_sc_hd__a21o_1 _19139_ (.A1(\rbzero.spi_registers.got_new_vinf ),
    .A2(_02724_),
    .B1(\rbzero.row_render.vinf ),
    .X(_02741_));
 sky130_fd_sc_hd__clkbuf_4 _19140_ (.A(_09243_),
    .X(_02742_));
 sky130_fd_sc_hd__o311a_1 _19141_ (.A1(\rbzero.spi_registers.new_vinf ),
    .A2(_02739_),
    .A3(_02740_),
    .B1(_02741_),
    .C1(_02742_),
    .X(_00742_));
 sky130_fd_sc_hd__and2_1 _19142_ (.A(\rbzero.spi_registers.got_new_leak ),
    .B(_02721_),
    .X(_02743_));
 sky130_fd_sc_hd__clkbuf_2 _19143_ (.A(_02743_),
    .X(_02744_));
 sky130_fd_sc_hd__nand2_1 _19144_ (.A(\rbzero.spi_registers.got_new_leak ),
    .B(_02724_),
    .Y(_02745_));
 sky130_fd_sc_hd__or2_1 _19145_ (.A(\rbzero.spi_registers.new_leak[0] ),
    .B(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__o211a_1 _19146_ (.A1(\rbzero.floor_leak[0] ),
    .A2(_02744_),
    .B1(_02746_),
    .C1(_02738_),
    .X(_00743_));
 sky130_fd_sc_hd__or2_1 _19147_ (.A(\rbzero.spi_registers.new_leak[1] ),
    .B(_02745_),
    .X(_02747_));
 sky130_fd_sc_hd__o211a_1 _19148_ (.A1(\rbzero.floor_leak[1] ),
    .A2(_02744_),
    .B1(_02747_),
    .C1(_02738_),
    .X(_00744_));
 sky130_fd_sc_hd__or2_1 _19149_ (.A(\rbzero.spi_registers.new_leak[2] ),
    .B(_02745_),
    .X(_02748_));
 sky130_fd_sc_hd__o211a_1 _19150_ (.A1(\rbzero.floor_leak[2] ),
    .A2(_02744_),
    .B1(_02748_),
    .C1(_02738_),
    .X(_00745_));
 sky130_fd_sc_hd__or2_1 _19151_ (.A(\rbzero.spi_registers.new_leak[3] ),
    .B(_02745_),
    .X(_02749_));
 sky130_fd_sc_hd__o211a_1 _19152_ (.A1(\rbzero.floor_leak[3] ),
    .A2(_02744_),
    .B1(_02749_),
    .C1(_02738_),
    .X(_00746_));
 sky130_fd_sc_hd__or2_1 _19153_ (.A(\rbzero.spi_registers.new_leak[4] ),
    .B(_02745_),
    .X(_02750_));
 sky130_fd_sc_hd__o211a_1 _19154_ (.A1(\rbzero.floor_leak[4] ),
    .A2(_02744_),
    .B1(_02750_),
    .C1(_02738_),
    .X(_00747_));
 sky130_fd_sc_hd__or2_1 _19155_ (.A(\rbzero.spi_registers.new_leak[5] ),
    .B(_02745_),
    .X(_02751_));
 sky130_fd_sc_hd__o211a_1 _19156_ (.A1(\rbzero.floor_leak[5] ),
    .A2(_02744_),
    .B1(_02751_),
    .C1(_02738_),
    .X(_00748_));
 sky130_fd_sc_hd__nand2_2 _19157_ (.A(\rbzero.spi_registers.got_new_sky ),
    .B(_02720_),
    .Y(_02752_));
 sky130_fd_sc_hd__buf_4 _19158_ (.A(_03442_),
    .X(_02753_));
 sky130_fd_sc_hd__a31o_1 _19159_ (.A1(\rbzero.spi_registers.new_sky[0] ),
    .A2(\rbzero.spi_registers.got_new_sky ),
    .A3(_02724_),
    .B1(_02753_),
    .X(_02754_));
 sky130_fd_sc_hd__a21o_1 _19160_ (.A1(\rbzero.color_sky[0] ),
    .A2(_02752_),
    .B1(_02754_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _19161_ (.A0(\rbzero.spi_registers.new_sky[1] ),
    .A1(\rbzero.color_sky[1] ),
    .S(_02752_),
    .X(_02755_));
 sky130_fd_sc_hd__and2_1 _19162_ (.A(_02742_),
    .B(_02755_),
    .X(_02756_));
 sky130_fd_sc_hd__clkbuf_1 _19163_ (.A(_02756_),
    .X(_00750_));
 sky130_fd_sc_hd__a31o_1 _19164_ (.A1(\rbzero.spi_registers.new_sky[2] ),
    .A2(\rbzero.spi_registers.got_new_sky ),
    .A3(_02724_),
    .B1(_02753_),
    .X(_02757_));
 sky130_fd_sc_hd__a21o_1 _19165_ (.A1(\rbzero.color_sky[2] ),
    .A2(_02752_),
    .B1(_02757_),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _19166_ (.A0(\rbzero.spi_registers.new_sky[3] ),
    .A1(\rbzero.color_sky[3] ),
    .S(_02752_),
    .X(_02758_));
 sky130_fd_sc_hd__and2_1 _19167_ (.A(_09247_),
    .B(_02758_),
    .X(_02759_));
 sky130_fd_sc_hd__clkbuf_1 _19168_ (.A(_02759_),
    .X(_00752_));
 sky130_fd_sc_hd__a31o_1 _19169_ (.A1(\rbzero.spi_registers.new_sky[4] ),
    .A2(\rbzero.spi_registers.got_new_sky ),
    .A3(_02724_),
    .B1(_02753_),
    .X(_02760_));
 sky130_fd_sc_hd__a21o_1 _19170_ (.A1(\rbzero.color_sky[4] ),
    .A2(_02752_),
    .B1(_02760_),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _19171_ (.A0(\rbzero.spi_registers.new_sky[5] ),
    .A1(\rbzero.color_sky[5] ),
    .S(_02752_),
    .X(_02761_));
 sky130_fd_sc_hd__and2_1 _19172_ (.A(_09247_),
    .B(_02761_),
    .X(_02762_));
 sky130_fd_sc_hd__clkbuf_1 _19173_ (.A(_02762_),
    .X(_00754_));
 sky130_fd_sc_hd__nand2_2 _19174_ (.A(\rbzero.spi_registers.got_new_floor ),
    .B(_02720_),
    .Y(_02763_));
 sky130_fd_sc_hd__mux2_1 _19175_ (.A0(\rbzero.spi_registers.new_floor[0] ),
    .A1(\rbzero.color_floor[0] ),
    .S(_02763_),
    .X(_02764_));
 sky130_fd_sc_hd__and2_1 _19176_ (.A(_09247_),
    .B(_02764_),
    .X(_02765_));
 sky130_fd_sc_hd__clkbuf_1 _19177_ (.A(_02765_),
    .X(_00755_));
 sky130_fd_sc_hd__a31o_1 _19178_ (.A1(\rbzero.spi_registers.new_floor[1] ),
    .A2(\rbzero.spi_registers.got_new_floor ),
    .A3(_02724_),
    .B1(_02753_),
    .X(_02766_));
 sky130_fd_sc_hd__a21o_1 _19179_ (.A1(\rbzero.color_floor[1] ),
    .A2(_02763_),
    .B1(_02766_),
    .X(_00756_));
 sky130_fd_sc_hd__mux2_1 _19180_ (.A0(\rbzero.spi_registers.new_floor[2] ),
    .A1(\rbzero.color_floor[2] ),
    .S(_02763_),
    .X(_02767_));
 sky130_fd_sc_hd__and2_1 _19181_ (.A(_09247_),
    .B(_02767_),
    .X(_02768_));
 sky130_fd_sc_hd__clkbuf_1 _19182_ (.A(_02768_),
    .X(_00757_));
 sky130_fd_sc_hd__a31o_1 _19183_ (.A1(\rbzero.spi_registers.new_floor[3] ),
    .A2(\rbzero.spi_registers.got_new_floor ),
    .A3(_02724_),
    .B1(_02753_),
    .X(_02769_));
 sky130_fd_sc_hd__a21o_1 _19184_ (.A1(\rbzero.color_floor[3] ),
    .A2(_02763_),
    .B1(_02769_),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_1 _19185_ (.A0(\rbzero.spi_registers.new_floor[4] ),
    .A1(\rbzero.color_floor[4] ),
    .S(_02763_),
    .X(_02770_));
 sky130_fd_sc_hd__and2_1 _19186_ (.A(_09247_),
    .B(_02770_),
    .X(_02771_));
 sky130_fd_sc_hd__clkbuf_1 _19187_ (.A(_02771_),
    .X(_00759_));
 sky130_fd_sc_hd__a31o_1 _19188_ (.A1(\rbzero.spi_registers.new_floor[5] ),
    .A2(\rbzero.spi_registers.got_new_floor ),
    .A3(_02724_),
    .B1(_02753_),
    .X(_02772_));
 sky130_fd_sc_hd__a21o_1 _19189_ (.A1(\rbzero.color_floor[5] ),
    .A2(_02763_),
    .B1(_02772_),
    .X(_00760_));
 sky130_fd_sc_hd__and2_1 _19190_ (.A(\rbzero.spi_registers.got_new_vshift ),
    .B(_02721_),
    .X(_02773_));
 sky130_fd_sc_hd__clkbuf_2 _19191_ (.A(_02773_),
    .X(_02774_));
 sky130_fd_sc_hd__nand2_1 _19192_ (.A(\rbzero.spi_registers.got_new_vshift ),
    .B(_02724_),
    .Y(_02775_));
 sky130_fd_sc_hd__or2_1 _19193_ (.A(\rbzero.spi_registers.new_vshift[0] ),
    .B(_02775_),
    .X(_02776_));
 sky130_fd_sc_hd__o211a_1 _19194_ (.A1(\rbzero.spi_registers.vshift[0] ),
    .A2(_02774_),
    .B1(_02776_),
    .C1(_02738_),
    .X(_00761_));
 sky130_fd_sc_hd__or2_1 _19195_ (.A(\rbzero.spi_registers.new_vshift[1] ),
    .B(_02775_),
    .X(_02777_));
 sky130_fd_sc_hd__o211a_1 _19196_ (.A1(\rbzero.spi_registers.vshift[1] ),
    .A2(_02774_),
    .B1(_02777_),
    .C1(_02738_),
    .X(_00762_));
 sky130_fd_sc_hd__or2_1 _19197_ (.A(\rbzero.spi_registers.new_vshift[2] ),
    .B(_02775_),
    .X(_02778_));
 sky130_fd_sc_hd__o211a_1 _19198_ (.A1(\rbzero.spi_registers.vshift[2] ),
    .A2(_02774_),
    .B1(_02778_),
    .C1(_02738_),
    .X(_00763_));
 sky130_fd_sc_hd__or2_1 _19199_ (.A(\rbzero.spi_registers.new_vshift[3] ),
    .B(_02775_),
    .X(_02779_));
 sky130_fd_sc_hd__buf_4 _19200_ (.A(_02727_),
    .X(_02780_));
 sky130_fd_sc_hd__o211a_1 _19201_ (.A1(\rbzero.spi_registers.vshift[3] ),
    .A2(_02774_),
    .B1(_02779_),
    .C1(_02780_),
    .X(_00764_));
 sky130_fd_sc_hd__or2_1 _19202_ (.A(\rbzero.spi_registers.new_vshift[4] ),
    .B(_02775_),
    .X(_02781_));
 sky130_fd_sc_hd__o211a_1 _19203_ (.A1(\rbzero.spi_registers.vshift[4] ),
    .A2(_02774_),
    .B1(_02781_),
    .C1(_02780_),
    .X(_00765_));
 sky130_fd_sc_hd__or2_1 _19204_ (.A(\rbzero.spi_registers.new_vshift[5] ),
    .B(_02775_),
    .X(_02782_));
 sky130_fd_sc_hd__o211a_1 _19205_ (.A1(\rbzero.spi_registers.vshift[5] ),
    .A2(_02774_),
    .B1(_02782_),
    .C1(_02780_),
    .X(_00766_));
 sky130_fd_sc_hd__and4b_1 _19206_ (.A_N(\rbzero.spi_registers.spi_done ),
    .B(_02589_),
    .C(_02576_),
    .D(_02587_),
    .X(_02783_));
 sky130_fd_sc_hd__clkbuf_1 _19207_ (.A(_02783_),
    .X(_00767_));
 sky130_fd_sc_hd__or4b_1 _19208_ (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .B(\rbzero.spi_registers.spi_cmd[2] ),
    .C(_03442_),
    .D_N(\rbzero.spi_registers.spi_done ),
    .X(_02784_));
 sky130_fd_sc_hd__or2_1 _19209_ (.A(_02578_),
    .B(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__clkbuf_4 _19210_ (.A(_02785_),
    .X(_02786_));
 sky130_fd_sc_hd__mux2_1 _19211_ (.A0(\rbzero.spi_registers.spi_buffer[0] ),
    .A1(\rbzero.spi_registers.new_sky[0] ),
    .S(_02786_),
    .X(_02787_));
 sky130_fd_sc_hd__clkbuf_1 _19212_ (.A(_02787_),
    .X(_00768_));
 sky130_fd_sc_hd__mux2_1 _19213_ (.A0(\rbzero.spi_registers.spi_buffer[1] ),
    .A1(\rbzero.spi_registers.new_sky[1] ),
    .S(_02786_),
    .X(_02788_));
 sky130_fd_sc_hd__clkbuf_1 _19214_ (.A(_02788_),
    .X(_00769_));
 sky130_fd_sc_hd__mux2_1 _19215_ (.A0(\rbzero.spi_registers.spi_buffer[2] ),
    .A1(\rbzero.spi_registers.new_sky[2] ),
    .S(_02786_),
    .X(_02789_));
 sky130_fd_sc_hd__clkbuf_1 _19216_ (.A(_02789_),
    .X(_00770_));
 sky130_fd_sc_hd__mux2_1 _19217_ (.A0(\rbzero.spi_registers.spi_buffer[3] ),
    .A1(\rbzero.spi_registers.new_sky[3] ),
    .S(_02786_),
    .X(_02790_));
 sky130_fd_sc_hd__clkbuf_1 _19218_ (.A(_02790_),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_1 _19219_ (.A0(\rbzero.spi_registers.spi_buffer[4] ),
    .A1(\rbzero.spi_registers.new_sky[4] ),
    .S(_02786_),
    .X(_02791_));
 sky130_fd_sc_hd__clkbuf_1 _19220_ (.A(_02791_),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _19221_ (.A0(\rbzero.spi_registers.spi_buffer[5] ),
    .A1(\rbzero.spi_registers.new_sky[5] ),
    .S(_02786_),
    .X(_02792_));
 sky130_fd_sc_hd__clkbuf_1 _19222_ (.A(_02792_),
    .X(_00773_));
 sky130_fd_sc_hd__inv_2 _19223_ (.A(_02786_),
    .Y(_02793_));
 sky130_fd_sc_hd__a31o_1 _19224_ (.A1(\rbzero.spi_registers.got_new_sky ),
    .A2(_02742_),
    .A3(_02740_),
    .B1(_02793_),
    .X(_00774_));
 sky130_fd_sc_hd__or3b_1 _19225_ (.A(_02784_),
    .B(\rbzero.spi_registers.spi_cmd[1] ),
    .C_N(\rbzero.spi_registers.spi_cmd[0] ),
    .X(_02794_));
 sky130_fd_sc_hd__clkbuf_4 _19226_ (.A(_02794_),
    .X(_02795_));
 sky130_fd_sc_hd__mux2_1 _19227_ (.A0(\rbzero.spi_registers.spi_buffer[0] ),
    .A1(\rbzero.spi_registers.new_floor[0] ),
    .S(_02795_),
    .X(_02796_));
 sky130_fd_sc_hd__clkbuf_1 _19228_ (.A(_02796_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _19229_ (.A0(\rbzero.spi_registers.spi_buffer[1] ),
    .A1(\rbzero.spi_registers.new_floor[1] ),
    .S(_02795_),
    .X(_02797_));
 sky130_fd_sc_hd__clkbuf_1 _19230_ (.A(_02797_),
    .X(_00776_));
 sky130_fd_sc_hd__mux2_1 _19231_ (.A0(\rbzero.spi_registers.spi_buffer[2] ),
    .A1(\rbzero.spi_registers.new_floor[2] ),
    .S(_02795_),
    .X(_02798_));
 sky130_fd_sc_hd__clkbuf_1 _19232_ (.A(_02798_),
    .X(_00777_));
 sky130_fd_sc_hd__mux2_1 _19233_ (.A0(\rbzero.spi_registers.spi_buffer[3] ),
    .A1(\rbzero.spi_registers.new_floor[3] ),
    .S(_02795_),
    .X(_02799_));
 sky130_fd_sc_hd__clkbuf_1 _19234_ (.A(_02799_),
    .X(_00778_));
 sky130_fd_sc_hd__mux2_1 _19235_ (.A0(\rbzero.spi_registers.spi_buffer[4] ),
    .A1(\rbzero.spi_registers.new_floor[4] ),
    .S(_02795_),
    .X(_02800_));
 sky130_fd_sc_hd__clkbuf_1 _19236_ (.A(_02800_),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_1 _19237_ (.A0(\rbzero.spi_registers.spi_buffer[5] ),
    .A1(\rbzero.spi_registers.new_floor[5] ),
    .S(_02795_),
    .X(_02801_));
 sky130_fd_sc_hd__clkbuf_1 _19238_ (.A(_02801_),
    .X(_00780_));
 sky130_fd_sc_hd__inv_2 _19239_ (.A(_02795_),
    .Y(_02802_));
 sky130_fd_sc_hd__a31o_1 _19240_ (.A1(\rbzero.spi_registers.got_new_floor ),
    .A2(_02742_),
    .A3(_02740_),
    .B1(_02802_),
    .X(_00781_));
 sky130_fd_sc_hd__or3b_1 _19241_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .B(_02784_),
    .C_N(\rbzero.spi_registers.spi_cmd[1] ),
    .X(_02803_));
 sky130_fd_sc_hd__buf_2 _19242_ (.A(_02803_),
    .X(_02804_));
 sky130_fd_sc_hd__mux2_1 _19243_ (.A0(\rbzero.spi_registers.spi_buffer[0] ),
    .A1(\rbzero.spi_registers.new_leak[0] ),
    .S(_02804_),
    .X(_02805_));
 sky130_fd_sc_hd__clkbuf_1 _19244_ (.A(_02805_),
    .X(_00782_));
 sky130_fd_sc_hd__mux2_1 _19245_ (.A0(\rbzero.spi_registers.spi_buffer[1] ),
    .A1(\rbzero.spi_registers.new_leak[1] ),
    .S(_02804_),
    .X(_02806_));
 sky130_fd_sc_hd__clkbuf_1 _19246_ (.A(_02806_),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _19247_ (.A0(\rbzero.spi_registers.spi_buffer[2] ),
    .A1(\rbzero.spi_registers.new_leak[2] ),
    .S(_02804_),
    .X(_02807_));
 sky130_fd_sc_hd__clkbuf_1 _19248_ (.A(_02807_),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _19249_ (.A0(\rbzero.spi_registers.spi_buffer[3] ),
    .A1(\rbzero.spi_registers.new_leak[3] ),
    .S(_02804_),
    .X(_02808_));
 sky130_fd_sc_hd__clkbuf_1 _19250_ (.A(_02808_),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _19251_ (.A0(\rbzero.spi_registers.spi_buffer[4] ),
    .A1(\rbzero.spi_registers.new_leak[4] ),
    .S(_02804_),
    .X(_02809_));
 sky130_fd_sc_hd__clkbuf_1 _19252_ (.A(_02809_),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _19253_ (.A0(\rbzero.spi_registers.spi_buffer[5] ),
    .A1(\rbzero.spi_registers.new_leak[5] ),
    .S(_02804_),
    .X(_02810_));
 sky130_fd_sc_hd__clkbuf_1 _19254_ (.A(_02810_),
    .X(_00787_));
 sky130_fd_sc_hd__inv_2 _19255_ (.A(_02804_),
    .Y(_02811_));
 sky130_fd_sc_hd__a31o_1 _19256_ (.A1(\rbzero.spi_registers.got_new_leak ),
    .A2(_02742_),
    .A3(_02740_),
    .B1(_02811_),
    .X(_00788_));
 sky130_fd_sc_hd__and3_1 _19257_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_03292_),
    .C(_02582_),
    .X(_02812_));
 sky130_fd_sc_hd__clkbuf_4 _19258_ (.A(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_1 _19259_ (.A0(\rbzero.spi_registers.new_other[0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__clkbuf_1 _19260_ (.A(_02814_),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _19261_ (.A0(\rbzero.spi_registers.new_other[1] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_02813_),
    .X(_02815_));
 sky130_fd_sc_hd__clkbuf_1 _19262_ (.A(_02815_),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _19263_ (.A0(\rbzero.spi_registers.new_other[2] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_02813_),
    .X(_02816_));
 sky130_fd_sc_hd__clkbuf_1 _19264_ (.A(_02816_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _19265_ (.A0(\rbzero.spi_registers.new_other[3] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_02813_),
    .X(_02817_));
 sky130_fd_sc_hd__clkbuf_1 _19266_ (.A(_02817_),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _19267_ (.A0(\rbzero.spi_registers.new_other[4] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_02813_),
    .X(_02818_));
 sky130_fd_sc_hd__clkbuf_1 _19268_ (.A(_02818_),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _19269_ (.A0(\rbzero.spi_registers.new_other[6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_02813_),
    .X(_02819_));
 sky130_fd_sc_hd__clkbuf_1 _19270_ (.A(_02819_),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _19271_ (.A0(\rbzero.spi_registers.new_other[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_02813_),
    .X(_02820_));
 sky130_fd_sc_hd__clkbuf_1 _19272_ (.A(_02820_),
    .X(_00795_));
 sky130_fd_sc_hd__mux2_1 _19273_ (.A0(\rbzero.spi_registers.new_other[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_02813_),
    .X(_02821_));
 sky130_fd_sc_hd__clkbuf_1 _19274_ (.A(_02821_),
    .X(_00796_));
 sky130_fd_sc_hd__mux2_1 _19275_ (.A0(\rbzero.spi_registers.new_other[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_02813_),
    .X(_02822_));
 sky130_fd_sc_hd__clkbuf_1 _19276_ (.A(_02822_),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _19277_ (.A0(\rbzero.spi_registers.new_other[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_02812_),
    .X(_02823_));
 sky130_fd_sc_hd__clkbuf_1 _19278_ (.A(_02823_),
    .X(_00798_));
 sky130_fd_sc_hd__a31o_1 _19279_ (.A1(\rbzero.spi_registers.got_new_other ),
    .A2(_02742_),
    .A3(_02740_),
    .B1(_02813_),
    .X(_00799_));
 sky130_fd_sc_hd__or4b_1 _19280_ (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .B(_02581_),
    .C(_02578_),
    .D_N(\rbzero.spi_registers.spi_done ),
    .X(_02824_));
 sky130_fd_sc_hd__nor2_4 _19281_ (.A(_03442_),
    .B(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__mux2_1 _19282_ (.A0(\rbzero.spi_registers.new_vshift[0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__clkbuf_1 _19283_ (.A(_02826_),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _19284_ (.A0(\rbzero.spi_registers.new_vshift[1] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_02825_),
    .X(_02827_));
 sky130_fd_sc_hd__clkbuf_1 _19285_ (.A(_02827_),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _19286_ (.A0(\rbzero.spi_registers.new_vshift[2] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_02825_),
    .X(_02828_));
 sky130_fd_sc_hd__clkbuf_1 _19287_ (.A(_02828_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _19288_ (.A0(\rbzero.spi_registers.new_vshift[3] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_02825_),
    .X(_02829_));
 sky130_fd_sc_hd__clkbuf_1 _19289_ (.A(_02829_),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _19290_ (.A0(\rbzero.spi_registers.new_vshift[4] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_02825_),
    .X(_02830_));
 sky130_fd_sc_hd__clkbuf_1 _19291_ (.A(_02830_),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _19292_ (.A0(\rbzero.spi_registers.new_vshift[5] ),
    .A1(\rbzero.spi_registers.spi_buffer[5] ),
    .S(_02825_),
    .X(_02831_));
 sky130_fd_sc_hd__clkbuf_1 _19293_ (.A(_02831_),
    .X(_00805_));
 sky130_fd_sc_hd__a31o_1 _19294_ (.A1(\rbzero.spi_registers.got_new_vshift ),
    .A2(_02742_),
    .A3(_02740_),
    .B1(_02825_),
    .X(_00806_));
 sky130_fd_sc_hd__clkbuf_4 _19295_ (.A(_04920_),
    .X(_02832_));
 sky130_fd_sc_hd__nor2_4 _19296_ (.A(net40),
    .B(net39),
    .Y(_02833_));
 sky130_fd_sc_hd__or2_1 _19297_ (.A(_02740_),
    .B(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__buf_2 _19298_ (.A(_02834_),
    .X(_02835_));
 sky130_fd_sc_hd__buf_2 _19299_ (.A(_02835_),
    .X(_02836_));
 sky130_fd_sc_hd__o211a_1 _19300_ (.A1(\rbzero.pov.spi_done ),
    .A2(\rbzero.pov.ready ),
    .B1(_02832_),
    .C1(_02836_),
    .X(_00807_));
 sky130_fd_sc_hd__nor2b_2 _19301_ (.A(\rbzero.pov.sclk_buffer[2] ),
    .B_N(\rbzero.pov.sclk_buffer[1] ),
    .Y(_02837_));
 sky130_fd_sc_hd__nor2_2 _19302_ (.A(\rbzero.pov.ss_buffer[1] ),
    .B(_03442_),
    .Y(_02838_));
 sky130_fd_sc_hd__o21ai_1 _19303_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_02837_),
    .B1(_02838_),
    .Y(_02839_));
 sky130_fd_sc_hd__a21oi_1 _19304_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_02837_),
    .B1(_02839_),
    .Y(_00808_));
 sky130_fd_sc_hd__and3_1 _19305_ (.A(\rbzero.pov.spi_counter[1] ),
    .B(\rbzero.pov.spi_counter[0] ),
    .C(_02837_),
    .X(_02840_));
 sky130_fd_sc_hd__a21o_1 _19306_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_02837_),
    .B1(\rbzero.pov.spi_counter[1] ),
    .X(_02841_));
 sky130_fd_sc_hd__and4bb_1 _19307_ (.A_N(\rbzero.pov.spi_counter[5] ),
    .B_N(\rbzero.pov.spi_counter[4] ),
    .C(\rbzero.pov.spi_counter[3] ),
    .D(\rbzero.pov.spi_counter[6] ),
    .X(_02842_));
 sky130_fd_sc_hd__and4bb_1 _19308_ (.A_N(\rbzero.pov.spi_counter[2] ),
    .B_N(\rbzero.pov.spi_counter[1] ),
    .C(\rbzero.pov.spi_counter[0] ),
    .D(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__a21boi_1 _19309_ (.A1(_02837_),
    .A2(_02843_),
    .B1_N(_02838_),
    .Y(_02844_));
 sky130_fd_sc_hd__and3b_1 _19310_ (.A_N(_02840_),
    .B(_02841_),
    .C(_02844_),
    .X(_02845_));
 sky130_fd_sc_hd__clkbuf_1 _19311_ (.A(_02845_),
    .X(_00809_));
 sky130_fd_sc_hd__and2_1 _19312_ (.A(\rbzero.pov.spi_counter[2] ),
    .B(_02840_),
    .X(_02846_));
 sky130_fd_sc_hd__o21ai_1 _19313_ (.A1(\rbzero.pov.spi_counter[2] ),
    .A2(_02840_),
    .B1(_02838_),
    .Y(_02847_));
 sky130_fd_sc_hd__nor2_1 _19314_ (.A(_02846_),
    .B(_02847_),
    .Y(_00810_));
 sky130_fd_sc_hd__nand2_1 _19315_ (.A(\rbzero.pov.spi_counter[3] ),
    .B(_02846_),
    .Y(_02848_));
 sky130_fd_sc_hd__o211a_1 _19316_ (.A1(\rbzero.pov.spi_counter[3] ),
    .A2(_02846_),
    .B1(_02848_),
    .C1(_02844_),
    .X(_00811_));
 sky130_fd_sc_hd__and3_1 _19317_ (.A(\rbzero.pov.spi_counter[4] ),
    .B(\rbzero.pov.spi_counter[3] ),
    .C(_02846_),
    .X(_02849_));
 sky130_fd_sc_hd__a31o_1 _19318_ (.A1(\rbzero.pov.spi_counter[3] ),
    .A2(\rbzero.pov.spi_counter[2] ),
    .A3(_02840_),
    .B1(\rbzero.pov.spi_counter[4] ),
    .X(_02850_));
 sky130_fd_sc_hd__and3b_1 _19319_ (.A_N(_02849_),
    .B(_02838_),
    .C(_02850_),
    .X(_02851_));
 sky130_fd_sc_hd__clkbuf_1 _19320_ (.A(_02851_),
    .X(_00812_));
 sky130_fd_sc_hd__and2_1 _19321_ (.A(\rbzero.pov.spi_counter[5] ),
    .B(_02849_),
    .X(_02852_));
 sky130_fd_sc_hd__o21ai_1 _19322_ (.A1(\rbzero.pov.spi_counter[5] ),
    .A2(_02849_),
    .B1(_02838_),
    .Y(_02853_));
 sky130_fd_sc_hd__nor2_1 _19323_ (.A(_02852_),
    .B(_02853_),
    .Y(_00813_));
 sky130_fd_sc_hd__a21boi_1 _19324_ (.A1(\rbzero.pov.spi_counter[6] ),
    .A2(_02852_),
    .B1_N(_02844_),
    .Y(_02854_));
 sky130_fd_sc_hd__o21a_1 _19325_ (.A1(\rbzero.pov.spi_counter[6] ),
    .A2(_02852_),
    .B1(_02854_),
    .X(_00814_));
 sky130_fd_sc_hd__buf_4 _19326_ (.A(_04702_),
    .X(_02855_));
 sky130_fd_sc_hd__buf_4 _19327_ (.A(_02855_),
    .X(_02856_));
 sky130_fd_sc_hd__clkinv_2 _19328_ (.A(_02856_),
    .Y(_00017_));
 sky130_fd_sc_hd__clkinv_2 _19329_ (.A(_02856_),
    .Y(_00018_));
 sky130_fd_sc_hd__clkinv_2 _19330_ (.A(_02856_),
    .Y(_00019_));
 sky130_fd_sc_hd__clkinv_2 _19331_ (.A(_02856_),
    .Y(_00020_));
 sky130_fd_sc_hd__clkinv_2 _19332_ (.A(_02856_),
    .Y(_00021_));
 sky130_fd_sc_hd__clkinv_2 _19333_ (.A(_02856_),
    .Y(_00022_));
 sky130_fd_sc_hd__clkinv_2 _19334_ (.A(_02856_),
    .Y(_00023_));
 sky130_fd_sc_hd__clkinv_2 _19335_ (.A(_02856_),
    .Y(_00024_));
 sky130_fd_sc_hd__clkinv_2 _19336_ (.A(_02856_),
    .Y(_00025_));
 sky130_fd_sc_hd__clkinv_2 _19337_ (.A(_02856_),
    .Y(_00026_));
 sky130_fd_sc_hd__buf_4 _19338_ (.A(_02855_),
    .X(_02857_));
 sky130_fd_sc_hd__clkinv_2 _19339_ (.A(_02857_),
    .Y(_00027_));
 sky130_fd_sc_hd__clkinv_2 _19340_ (.A(_02857_),
    .Y(_00028_));
 sky130_fd_sc_hd__clkinv_2 _19341_ (.A(_02857_),
    .Y(_00029_));
 sky130_fd_sc_hd__clkinv_2 _19342_ (.A(_02857_),
    .Y(_00030_));
 sky130_fd_sc_hd__clkinv_2 _19343_ (.A(_02857_),
    .Y(_00031_));
 sky130_fd_sc_hd__clkinv_2 _19344_ (.A(_02857_),
    .Y(_00032_));
 sky130_fd_sc_hd__clkinv_2 _19345_ (.A(_02857_),
    .Y(_00033_));
 sky130_fd_sc_hd__clkinv_2 _19346_ (.A(_02857_),
    .Y(_00034_));
 sky130_fd_sc_hd__clkinv_2 _19347_ (.A(_02857_),
    .Y(_00035_));
 sky130_fd_sc_hd__clkinv_2 _19348_ (.A(_02857_),
    .Y(_00036_));
 sky130_fd_sc_hd__buf_4 _19349_ (.A(_02855_),
    .X(_02858_));
 sky130_fd_sc_hd__clkinv_2 _19350_ (.A(_02858_),
    .Y(_00037_));
 sky130_fd_sc_hd__clkinv_2 _19351_ (.A(_02858_),
    .Y(_00038_));
 sky130_fd_sc_hd__clkinv_2 _19352_ (.A(_02858_),
    .Y(_00039_));
 sky130_fd_sc_hd__clkinv_2 _19353_ (.A(_02858_),
    .Y(_00040_));
 sky130_fd_sc_hd__clkinv_2 _19354_ (.A(_02858_),
    .Y(_00041_));
 sky130_fd_sc_hd__clkinv_2 _19355_ (.A(_02858_),
    .Y(_00042_));
 sky130_fd_sc_hd__clkinv_2 _19356_ (.A(_02858_),
    .Y(_00043_));
 sky130_fd_sc_hd__clkinv_2 _19357_ (.A(_02858_),
    .Y(_00044_));
 sky130_fd_sc_hd__clkinv_2 _19358_ (.A(_02858_),
    .Y(_00045_));
 sky130_fd_sc_hd__clkinv_2 _19359_ (.A(_02858_),
    .Y(_00046_));
 sky130_fd_sc_hd__buf_4 _19360_ (.A(_02855_),
    .X(_02859_));
 sky130_fd_sc_hd__clkinv_2 _19361_ (.A(_02859_),
    .Y(_00047_));
 sky130_fd_sc_hd__clkinv_2 _19362_ (.A(_02859_),
    .Y(_00048_));
 sky130_fd_sc_hd__clkinv_2 _19363_ (.A(_02859_),
    .Y(_00049_));
 sky130_fd_sc_hd__clkinv_2 _19364_ (.A(_02859_),
    .Y(_00050_));
 sky130_fd_sc_hd__clkinv_2 _19365_ (.A(_02859_),
    .Y(_00051_));
 sky130_fd_sc_hd__clkinv_2 _19366_ (.A(_02859_),
    .Y(_00052_));
 sky130_fd_sc_hd__clkinv_2 _19367_ (.A(_02859_),
    .Y(_00053_));
 sky130_fd_sc_hd__clkinv_2 _19368_ (.A(_02859_),
    .Y(_00054_));
 sky130_fd_sc_hd__clkinv_2 _19369_ (.A(_02859_),
    .Y(_00055_));
 sky130_fd_sc_hd__clkinv_2 _19370_ (.A(_02859_),
    .Y(_00056_));
 sky130_fd_sc_hd__buf_4 _19371_ (.A(_02855_),
    .X(_02860_));
 sky130_fd_sc_hd__clkinv_2 _19372_ (.A(_02860_),
    .Y(_00057_));
 sky130_fd_sc_hd__clkinv_2 _19373_ (.A(_02860_),
    .Y(_00058_));
 sky130_fd_sc_hd__clkinv_2 _19374_ (.A(_02860_),
    .Y(_00059_));
 sky130_fd_sc_hd__clkinv_2 _19375_ (.A(_02860_),
    .Y(_00060_));
 sky130_fd_sc_hd__clkinv_2 _19376_ (.A(_02860_),
    .Y(_00061_));
 sky130_fd_sc_hd__clkinv_2 _19377_ (.A(_02860_),
    .Y(_00062_));
 sky130_fd_sc_hd__clkinv_2 _19378_ (.A(_02860_),
    .Y(_00063_));
 sky130_fd_sc_hd__clkinv_2 _19379_ (.A(_02860_),
    .Y(_00064_));
 sky130_fd_sc_hd__clkinv_2 _19380_ (.A(_02860_),
    .Y(_00065_));
 sky130_fd_sc_hd__clkinv_2 _19381_ (.A(_02860_),
    .Y(_00066_));
 sky130_fd_sc_hd__buf_4 _19382_ (.A(_02855_),
    .X(_02861_));
 sky130_fd_sc_hd__clkinv_2 _19383_ (.A(_02861_),
    .Y(_00067_));
 sky130_fd_sc_hd__clkinv_2 _19384_ (.A(_02861_),
    .Y(_00068_));
 sky130_fd_sc_hd__clkinv_2 _19385_ (.A(_02861_),
    .Y(_00069_));
 sky130_fd_sc_hd__clkinv_2 _19386_ (.A(_02861_),
    .Y(_00070_));
 sky130_fd_sc_hd__clkinv_2 _19387_ (.A(_02861_),
    .Y(_00071_));
 sky130_fd_sc_hd__clkinv_2 _19388_ (.A(_02861_),
    .Y(_00072_));
 sky130_fd_sc_hd__clkinv_2 _19389_ (.A(_02861_),
    .Y(_00073_));
 sky130_fd_sc_hd__clkinv_2 _19390_ (.A(_02861_),
    .Y(_00074_));
 sky130_fd_sc_hd__clkinv_2 _19391_ (.A(_02861_),
    .Y(_00075_));
 sky130_fd_sc_hd__clkinv_2 _19392_ (.A(_02861_),
    .Y(_00076_));
 sky130_fd_sc_hd__buf_4 _19393_ (.A(_04702_),
    .X(_02862_));
 sky130_fd_sc_hd__buf_4 _19394_ (.A(_02862_),
    .X(_02863_));
 sky130_fd_sc_hd__clkinv_2 _19395_ (.A(_02863_),
    .Y(_00077_));
 sky130_fd_sc_hd__clkinv_2 _19396_ (.A(_02863_),
    .Y(_00078_));
 sky130_fd_sc_hd__clkinv_2 _19397_ (.A(_02863_),
    .Y(_00079_));
 sky130_fd_sc_hd__clkinv_2 _19398_ (.A(_02863_),
    .Y(_00080_));
 sky130_fd_sc_hd__nand2_2 _19399_ (.A(_02838_),
    .B(_02837_),
    .Y(_02864_));
 sky130_fd_sc_hd__clkbuf_4 _19400_ (.A(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__clkbuf_4 _19401_ (.A(_02865_),
    .X(_02866_));
 sky130_fd_sc_hd__mux2_1 _19402_ (.A0(\rbzero.pov.mosi ),
    .A1(\rbzero.pov.spi_buffer[0] ),
    .S(_02866_),
    .X(_02867_));
 sky130_fd_sc_hd__clkbuf_1 _19403_ (.A(_02867_),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _19404_ (.A0(\rbzero.pov.spi_buffer[0] ),
    .A1(\rbzero.pov.spi_buffer[1] ),
    .S(_02866_),
    .X(_02868_));
 sky130_fd_sc_hd__clkbuf_1 _19405_ (.A(_02868_),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _19406_ (.A0(\rbzero.pov.spi_buffer[1] ),
    .A1(\rbzero.pov.spi_buffer[2] ),
    .S(_02866_),
    .X(_02869_));
 sky130_fd_sc_hd__clkbuf_1 _19407_ (.A(_02869_),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _19408_ (.A0(\rbzero.pov.spi_buffer[2] ),
    .A1(\rbzero.pov.spi_buffer[3] ),
    .S(_02866_),
    .X(_02870_));
 sky130_fd_sc_hd__clkbuf_1 _19409_ (.A(_02870_),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_1 _19410_ (.A0(\rbzero.pov.spi_buffer[3] ),
    .A1(\rbzero.pov.spi_buffer[4] ),
    .S(_02866_),
    .X(_02871_));
 sky130_fd_sc_hd__clkbuf_1 _19411_ (.A(_02871_),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_1 _19412_ (.A0(\rbzero.pov.spi_buffer[4] ),
    .A1(\rbzero.pov.spi_buffer[5] ),
    .S(_02866_),
    .X(_02872_));
 sky130_fd_sc_hd__clkbuf_1 _19413_ (.A(_02872_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _19414_ (.A0(\rbzero.pov.spi_buffer[5] ),
    .A1(\rbzero.pov.spi_buffer[6] ),
    .S(_02866_),
    .X(_02873_));
 sky130_fd_sc_hd__clkbuf_1 _19415_ (.A(_02873_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _19416_ (.A0(\rbzero.pov.spi_buffer[6] ),
    .A1(\rbzero.pov.spi_buffer[7] ),
    .S(_02866_),
    .X(_02874_));
 sky130_fd_sc_hd__clkbuf_1 _19417_ (.A(_02874_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _19418_ (.A0(\rbzero.pov.spi_buffer[7] ),
    .A1(\rbzero.pov.spi_buffer[8] ),
    .S(_02866_),
    .X(_02875_));
 sky130_fd_sc_hd__clkbuf_1 _19419_ (.A(_02875_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _19420_ (.A0(\rbzero.pov.spi_buffer[8] ),
    .A1(\rbzero.pov.spi_buffer[9] ),
    .S(_02866_),
    .X(_02876_));
 sky130_fd_sc_hd__clkbuf_1 _19421_ (.A(_02876_),
    .X(_00888_));
 sky130_fd_sc_hd__clkbuf_4 _19422_ (.A(_02865_),
    .X(_02877_));
 sky130_fd_sc_hd__mux2_1 _19423_ (.A0(\rbzero.pov.spi_buffer[9] ),
    .A1(\rbzero.pov.spi_buffer[10] ),
    .S(_02877_),
    .X(_02878_));
 sky130_fd_sc_hd__clkbuf_1 _19424_ (.A(_02878_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _19425_ (.A0(\rbzero.pov.spi_buffer[10] ),
    .A1(\rbzero.pov.spi_buffer[11] ),
    .S(_02877_),
    .X(_02879_));
 sky130_fd_sc_hd__clkbuf_1 _19426_ (.A(_02879_),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _19427_ (.A0(\rbzero.pov.spi_buffer[11] ),
    .A1(\rbzero.pov.spi_buffer[12] ),
    .S(_02877_),
    .X(_02880_));
 sky130_fd_sc_hd__clkbuf_1 _19428_ (.A(_02880_),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _19429_ (.A0(\rbzero.pov.spi_buffer[12] ),
    .A1(\rbzero.pov.spi_buffer[13] ),
    .S(_02877_),
    .X(_02881_));
 sky130_fd_sc_hd__clkbuf_1 _19430_ (.A(_02881_),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _19431_ (.A0(\rbzero.pov.spi_buffer[13] ),
    .A1(\rbzero.pov.spi_buffer[14] ),
    .S(_02877_),
    .X(_02882_));
 sky130_fd_sc_hd__clkbuf_1 _19432_ (.A(_02882_),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _19433_ (.A0(\rbzero.pov.spi_buffer[14] ),
    .A1(\rbzero.pov.spi_buffer[15] ),
    .S(_02877_),
    .X(_02883_));
 sky130_fd_sc_hd__clkbuf_1 _19434_ (.A(_02883_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _19435_ (.A0(\rbzero.pov.spi_buffer[15] ),
    .A1(\rbzero.pov.spi_buffer[16] ),
    .S(_02877_),
    .X(_02884_));
 sky130_fd_sc_hd__clkbuf_1 _19436_ (.A(_02884_),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_1 _19437_ (.A0(\rbzero.pov.spi_buffer[16] ),
    .A1(\rbzero.pov.spi_buffer[17] ),
    .S(_02877_),
    .X(_02885_));
 sky130_fd_sc_hd__clkbuf_1 _19438_ (.A(_02885_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _19439_ (.A0(\rbzero.pov.spi_buffer[17] ),
    .A1(\rbzero.pov.spi_buffer[18] ),
    .S(_02877_),
    .X(_02886_));
 sky130_fd_sc_hd__clkbuf_1 _19440_ (.A(_02886_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _19441_ (.A0(\rbzero.pov.spi_buffer[18] ),
    .A1(\rbzero.pov.spi_buffer[19] ),
    .S(_02877_),
    .X(_02887_));
 sky130_fd_sc_hd__clkbuf_1 _19442_ (.A(_02887_),
    .X(_00898_));
 sky130_fd_sc_hd__clkbuf_4 _19443_ (.A(_02865_),
    .X(_02888_));
 sky130_fd_sc_hd__mux2_1 _19444_ (.A0(\rbzero.pov.spi_buffer[19] ),
    .A1(\rbzero.pov.spi_buffer[20] ),
    .S(_02888_),
    .X(_02889_));
 sky130_fd_sc_hd__clkbuf_1 _19445_ (.A(_02889_),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _19446_ (.A0(\rbzero.pov.spi_buffer[20] ),
    .A1(\rbzero.pov.spi_buffer[21] ),
    .S(_02888_),
    .X(_02890_));
 sky130_fd_sc_hd__clkbuf_1 _19447_ (.A(_02890_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _19448_ (.A0(\rbzero.pov.spi_buffer[21] ),
    .A1(\rbzero.pov.spi_buffer[22] ),
    .S(_02888_),
    .X(_02891_));
 sky130_fd_sc_hd__clkbuf_1 _19449_ (.A(_02891_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _19450_ (.A0(\rbzero.pov.spi_buffer[22] ),
    .A1(\rbzero.pov.spi_buffer[23] ),
    .S(_02888_),
    .X(_02892_));
 sky130_fd_sc_hd__clkbuf_1 _19451_ (.A(_02892_),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _19452_ (.A0(\rbzero.pov.spi_buffer[23] ),
    .A1(\rbzero.pov.spi_buffer[24] ),
    .S(_02888_),
    .X(_02893_));
 sky130_fd_sc_hd__clkbuf_1 _19453_ (.A(_02893_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _19454_ (.A0(\rbzero.pov.spi_buffer[24] ),
    .A1(\rbzero.pov.spi_buffer[25] ),
    .S(_02888_),
    .X(_02894_));
 sky130_fd_sc_hd__clkbuf_1 _19455_ (.A(_02894_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _19456_ (.A0(\rbzero.pov.spi_buffer[25] ),
    .A1(\rbzero.pov.spi_buffer[26] ),
    .S(_02888_),
    .X(_02895_));
 sky130_fd_sc_hd__clkbuf_1 _19457_ (.A(_02895_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _19458_ (.A0(\rbzero.pov.spi_buffer[26] ),
    .A1(\rbzero.pov.spi_buffer[27] ),
    .S(_02888_),
    .X(_02896_));
 sky130_fd_sc_hd__clkbuf_1 _19459_ (.A(_02896_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _19460_ (.A0(\rbzero.pov.spi_buffer[27] ),
    .A1(\rbzero.pov.spi_buffer[28] ),
    .S(_02888_),
    .X(_02897_));
 sky130_fd_sc_hd__clkbuf_1 _19461_ (.A(_02897_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _19462_ (.A0(\rbzero.pov.spi_buffer[28] ),
    .A1(\rbzero.pov.spi_buffer[29] ),
    .S(_02888_),
    .X(_02898_));
 sky130_fd_sc_hd__clkbuf_1 _19463_ (.A(_02898_),
    .X(_00908_));
 sky130_fd_sc_hd__clkbuf_4 _19464_ (.A(_02865_),
    .X(_02899_));
 sky130_fd_sc_hd__mux2_1 _19465_ (.A0(\rbzero.pov.spi_buffer[29] ),
    .A1(\rbzero.pov.spi_buffer[30] ),
    .S(_02899_),
    .X(_02900_));
 sky130_fd_sc_hd__clkbuf_1 _19466_ (.A(_02900_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _19467_ (.A0(\rbzero.pov.spi_buffer[30] ),
    .A1(\rbzero.pov.spi_buffer[31] ),
    .S(_02899_),
    .X(_02901_));
 sky130_fd_sc_hd__clkbuf_1 _19468_ (.A(_02901_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _19469_ (.A0(\rbzero.pov.spi_buffer[31] ),
    .A1(\rbzero.pov.spi_buffer[32] ),
    .S(_02899_),
    .X(_02902_));
 sky130_fd_sc_hd__clkbuf_1 _19470_ (.A(_02902_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _19471_ (.A0(\rbzero.pov.spi_buffer[32] ),
    .A1(\rbzero.pov.spi_buffer[33] ),
    .S(_02899_),
    .X(_02903_));
 sky130_fd_sc_hd__clkbuf_1 _19472_ (.A(_02903_),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _19473_ (.A0(\rbzero.pov.spi_buffer[33] ),
    .A1(\rbzero.pov.spi_buffer[34] ),
    .S(_02899_),
    .X(_02904_));
 sky130_fd_sc_hd__clkbuf_1 _19474_ (.A(_02904_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _19475_ (.A0(\rbzero.pov.spi_buffer[34] ),
    .A1(\rbzero.pov.spi_buffer[35] ),
    .S(_02899_),
    .X(_02905_));
 sky130_fd_sc_hd__clkbuf_1 _19476_ (.A(_02905_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _19477_ (.A0(\rbzero.pov.spi_buffer[35] ),
    .A1(\rbzero.pov.spi_buffer[36] ),
    .S(_02899_),
    .X(_02906_));
 sky130_fd_sc_hd__clkbuf_1 _19478_ (.A(_02906_),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _19479_ (.A0(\rbzero.pov.spi_buffer[36] ),
    .A1(\rbzero.pov.spi_buffer[37] ),
    .S(_02899_),
    .X(_02907_));
 sky130_fd_sc_hd__clkbuf_1 _19480_ (.A(_02907_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _19481_ (.A0(\rbzero.pov.spi_buffer[37] ),
    .A1(\rbzero.pov.spi_buffer[38] ),
    .S(_02899_),
    .X(_02908_));
 sky130_fd_sc_hd__clkbuf_1 _19482_ (.A(_02908_),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _19483_ (.A0(\rbzero.pov.spi_buffer[38] ),
    .A1(\rbzero.pov.spi_buffer[39] ),
    .S(_02899_),
    .X(_02909_));
 sky130_fd_sc_hd__clkbuf_1 _19484_ (.A(_02909_),
    .X(_00918_));
 sky130_fd_sc_hd__clkbuf_4 _19485_ (.A(_02865_),
    .X(_02910_));
 sky130_fd_sc_hd__mux2_1 _19486_ (.A0(\rbzero.pov.spi_buffer[39] ),
    .A1(\rbzero.pov.spi_buffer[40] ),
    .S(_02910_),
    .X(_02911_));
 sky130_fd_sc_hd__clkbuf_1 _19487_ (.A(_02911_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _19488_ (.A0(\rbzero.pov.spi_buffer[40] ),
    .A1(\rbzero.pov.spi_buffer[41] ),
    .S(_02910_),
    .X(_02912_));
 sky130_fd_sc_hd__clkbuf_1 _19489_ (.A(_02912_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _19490_ (.A0(\rbzero.pov.spi_buffer[41] ),
    .A1(\rbzero.pov.spi_buffer[42] ),
    .S(_02910_),
    .X(_02913_));
 sky130_fd_sc_hd__clkbuf_1 _19491_ (.A(_02913_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _19492_ (.A0(\rbzero.pov.spi_buffer[42] ),
    .A1(\rbzero.pov.spi_buffer[43] ),
    .S(_02910_),
    .X(_02914_));
 sky130_fd_sc_hd__clkbuf_1 _19493_ (.A(_02914_),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _19494_ (.A0(\rbzero.pov.spi_buffer[43] ),
    .A1(\rbzero.pov.spi_buffer[44] ),
    .S(_02910_),
    .X(_02915_));
 sky130_fd_sc_hd__clkbuf_1 _19495_ (.A(_02915_),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_1 _19496_ (.A0(\rbzero.pov.spi_buffer[44] ),
    .A1(\rbzero.pov.spi_buffer[45] ),
    .S(_02910_),
    .X(_02916_));
 sky130_fd_sc_hd__clkbuf_1 _19497_ (.A(_02916_),
    .X(_00924_));
 sky130_fd_sc_hd__mux2_1 _19498_ (.A0(\rbzero.pov.spi_buffer[45] ),
    .A1(\rbzero.pov.spi_buffer[46] ),
    .S(_02910_),
    .X(_02917_));
 sky130_fd_sc_hd__clkbuf_1 _19499_ (.A(_02917_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _19500_ (.A0(\rbzero.pov.spi_buffer[46] ),
    .A1(\rbzero.pov.spi_buffer[47] ),
    .S(_02910_),
    .X(_02918_));
 sky130_fd_sc_hd__clkbuf_1 _19501_ (.A(_02918_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _19502_ (.A0(\rbzero.pov.spi_buffer[47] ),
    .A1(\rbzero.pov.spi_buffer[48] ),
    .S(_02910_),
    .X(_02919_));
 sky130_fd_sc_hd__clkbuf_1 _19503_ (.A(_02919_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _19504_ (.A0(\rbzero.pov.spi_buffer[48] ),
    .A1(\rbzero.pov.spi_buffer[49] ),
    .S(_02910_),
    .X(_02920_));
 sky130_fd_sc_hd__clkbuf_1 _19505_ (.A(_02920_),
    .X(_00928_));
 sky130_fd_sc_hd__clkbuf_4 _19506_ (.A(_02865_),
    .X(_02921_));
 sky130_fd_sc_hd__mux2_1 _19507_ (.A0(\rbzero.pov.spi_buffer[49] ),
    .A1(\rbzero.pov.spi_buffer[50] ),
    .S(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__clkbuf_1 _19508_ (.A(_02922_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _19509_ (.A0(\rbzero.pov.spi_buffer[50] ),
    .A1(\rbzero.pov.spi_buffer[51] ),
    .S(_02921_),
    .X(_02923_));
 sky130_fd_sc_hd__clkbuf_1 _19510_ (.A(_02923_),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _19511_ (.A0(\rbzero.pov.spi_buffer[51] ),
    .A1(\rbzero.pov.spi_buffer[52] ),
    .S(_02921_),
    .X(_02924_));
 sky130_fd_sc_hd__clkbuf_1 _19512_ (.A(_02924_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _19513_ (.A0(\rbzero.pov.spi_buffer[52] ),
    .A1(\rbzero.pov.spi_buffer[53] ),
    .S(_02921_),
    .X(_02925_));
 sky130_fd_sc_hd__clkbuf_1 _19514_ (.A(_02925_),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _19515_ (.A0(\rbzero.pov.spi_buffer[53] ),
    .A1(\rbzero.pov.spi_buffer[54] ),
    .S(_02921_),
    .X(_02926_));
 sky130_fd_sc_hd__clkbuf_1 _19516_ (.A(_02926_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _19517_ (.A0(\rbzero.pov.spi_buffer[54] ),
    .A1(\rbzero.pov.spi_buffer[55] ),
    .S(_02921_),
    .X(_02927_));
 sky130_fd_sc_hd__clkbuf_1 _19518_ (.A(_02927_),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _19519_ (.A0(\rbzero.pov.spi_buffer[55] ),
    .A1(\rbzero.pov.spi_buffer[56] ),
    .S(_02921_),
    .X(_02928_));
 sky130_fd_sc_hd__clkbuf_1 _19520_ (.A(_02928_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _19521_ (.A0(\rbzero.pov.spi_buffer[56] ),
    .A1(\rbzero.pov.spi_buffer[57] ),
    .S(_02921_),
    .X(_02929_));
 sky130_fd_sc_hd__clkbuf_1 _19522_ (.A(_02929_),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _19523_ (.A0(\rbzero.pov.spi_buffer[57] ),
    .A1(\rbzero.pov.spi_buffer[58] ),
    .S(_02921_),
    .X(_02930_));
 sky130_fd_sc_hd__clkbuf_1 _19524_ (.A(_02930_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _19525_ (.A0(\rbzero.pov.spi_buffer[58] ),
    .A1(\rbzero.pov.spi_buffer[59] ),
    .S(_02921_),
    .X(_02931_));
 sky130_fd_sc_hd__clkbuf_1 _19526_ (.A(_02931_),
    .X(_00938_));
 sky130_fd_sc_hd__clkbuf_4 _19527_ (.A(_02864_),
    .X(_02932_));
 sky130_fd_sc_hd__mux2_1 _19528_ (.A0(\rbzero.pov.spi_buffer[59] ),
    .A1(\rbzero.pov.spi_buffer[60] ),
    .S(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__clkbuf_1 _19529_ (.A(_02933_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _19530_ (.A0(\rbzero.pov.spi_buffer[60] ),
    .A1(\rbzero.pov.spi_buffer[61] ),
    .S(_02932_),
    .X(_02934_));
 sky130_fd_sc_hd__clkbuf_1 _19531_ (.A(_02934_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _19532_ (.A0(\rbzero.pov.spi_buffer[61] ),
    .A1(\rbzero.pov.spi_buffer[62] ),
    .S(_02932_),
    .X(_02935_));
 sky130_fd_sc_hd__clkbuf_1 _19533_ (.A(_02935_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _19534_ (.A0(\rbzero.pov.spi_buffer[62] ),
    .A1(\rbzero.pov.spi_buffer[63] ),
    .S(_02932_),
    .X(_02936_));
 sky130_fd_sc_hd__clkbuf_1 _19535_ (.A(_02936_),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _19536_ (.A0(\rbzero.pov.spi_buffer[63] ),
    .A1(\rbzero.pov.spi_buffer[64] ),
    .S(_02932_),
    .X(_02937_));
 sky130_fd_sc_hd__clkbuf_1 _19537_ (.A(_02937_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _19538_ (.A0(\rbzero.pov.spi_buffer[64] ),
    .A1(\rbzero.pov.spi_buffer[65] ),
    .S(_02932_),
    .X(_02938_));
 sky130_fd_sc_hd__clkbuf_1 _19539_ (.A(_02938_),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _19540_ (.A0(\rbzero.pov.spi_buffer[65] ),
    .A1(\rbzero.pov.spi_buffer[66] ),
    .S(_02932_),
    .X(_02939_));
 sky130_fd_sc_hd__clkbuf_1 _19541_ (.A(_02939_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _19542_ (.A0(\rbzero.pov.spi_buffer[66] ),
    .A1(\rbzero.pov.spi_buffer[67] ),
    .S(_02932_),
    .X(_02940_));
 sky130_fd_sc_hd__clkbuf_1 _19543_ (.A(_02940_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _19544_ (.A0(\rbzero.pov.spi_buffer[67] ),
    .A1(\rbzero.pov.spi_buffer[68] ),
    .S(_02932_),
    .X(_02941_));
 sky130_fd_sc_hd__clkbuf_1 _19545_ (.A(_02941_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _19546_ (.A0(\rbzero.pov.spi_buffer[68] ),
    .A1(\rbzero.pov.spi_buffer[69] ),
    .S(_02932_),
    .X(_02942_));
 sky130_fd_sc_hd__clkbuf_1 _19547_ (.A(_02942_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _19548_ (.A0(\rbzero.pov.spi_buffer[69] ),
    .A1(\rbzero.pov.spi_buffer[70] ),
    .S(_02865_),
    .X(_02943_));
 sky130_fd_sc_hd__clkbuf_1 _19549_ (.A(_02943_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _19550_ (.A0(\rbzero.pov.spi_buffer[70] ),
    .A1(\rbzero.pov.spi_buffer[71] ),
    .S(_02865_),
    .X(_02944_));
 sky130_fd_sc_hd__clkbuf_1 _19551_ (.A(_02944_),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _19552_ (.A0(\rbzero.pov.spi_buffer[71] ),
    .A1(\rbzero.pov.spi_buffer[72] ),
    .S(_02865_),
    .X(_02945_));
 sky130_fd_sc_hd__clkbuf_1 _19553_ (.A(_02945_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _19554_ (.A0(\rbzero.pov.spi_buffer[72] ),
    .A1(\rbzero.pov.spi_buffer[73] ),
    .S(_02865_),
    .X(_02946_));
 sky130_fd_sc_hd__clkbuf_1 _19555_ (.A(_02946_),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _19556_ (.A0(net52),
    .A1(\rbzero.pov.mosi_buffer[0] ),
    .S(_02708_),
    .X(_02947_));
 sky130_fd_sc_hd__clkbuf_1 _19557_ (.A(_02947_),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _19558_ (.A0(\rbzero.pov.mosi ),
    .A1(\rbzero.pov.mosi_buffer[0] ),
    .S(_09243_),
    .X(_02948_));
 sky130_fd_sc_hd__clkbuf_1 _19559_ (.A(_02948_),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _19560_ (.A0(net51),
    .A1(\rbzero.pov.ss_buffer[0] ),
    .S(_02708_),
    .X(_02949_));
 sky130_fd_sc_hd__clkbuf_1 _19561_ (.A(_02949_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _19562_ (.A0(\rbzero.pov.ss_buffer[1] ),
    .A1(\rbzero.pov.ss_buffer[0] ),
    .S(_09243_),
    .X(_02950_));
 sky130_fd_sc_hd__clkbuf_1 _19563_ (.A(_02950_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _19564_ (.A0(net53),
    .A1(\rbzero.pov.sclk_buffer[0] ),
    .S(_02708_),
    .X(_02951_));
 sky130_fd_sc_hd__clkbuf_1 _19565_ (.A(_02951_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _19566_ (.A0(\rbzero.pov.sclk_buffer[1] ),
    .A1(\rbzero.pov.sclk_buffer[0] ),
    .S(_09243_),
    .X(_02952_));
 sky130_fd_sc_hd__clkbuf_1 _19567_ (.A(_02952_),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _19568_ (.A0(\rbzero.pov.sclk_buffer[2] ),
    .A1(\rbzero.pov.sclk_buffer[1] ),
    .S(_09243_),
    .X(_02953_));
 sky130_fd_sc_hd__clkbuf_1 _19569_ (.A(_02953_),
    .X(_00959_));
 sky130_fd_sc_hd__and2_2 _19570_ (.A(\rbzero.pov.ready ),
    .B(_02834_),
    .X(_02954_));
 sky130_fd_sc_hd__o21ai_4 _19571_ (.A1(net39),
    .A2(_02954_),
    .B1(_02721_),
    .Y(_02955_));
 sky130_fd_sc_hd__clkbuf_4 _19572_ (.A(_02955_),
    .X(_02956_));
 sky130_fd_sc_hd__inv_2 _19573_ (.A(\rbzero.debug_overlay.playerX[-9] ),
    .Y(_02957_));
 sky130_fd_sc_hd__buf_2 _19574_ (.A(_02834_),
    .X(_02958_));
 sky130_fd_sc_hd__mux2_1 _19575_ (.A0(_02957_),
    .A1(\rbzero.pov.ready_buffer[59] ),
    .S(_02958_),
    .X(_02959_));
 sky130_fd_sc_hd__clkbuf_4 _19576_ (.A(_02955_),
    .X(_02960_));
 sky130_fd_sc_hd__nand2_1 _19577_ (.A(_02957_),
    .B(_02960_),
    .Y(_02961_));
 sky130_fd_sc_hd__o211a_1 _19578_ (.A1(_02956_),
    .A2(_02959_),
    .B1(_02961_),
    .C1(_02780_),
    .X(_00960_));
 sky130_fd_sc_hd__nor2_4 _19579_ (.A(_02740_),
    .B(_02833_),
    .Y(_02962_));
 sky130_fd_sc_hd__clkbuf_4 _19580_ (.A(_02962_),
    .X(_02963_));
 sky130_fd_sc_hd__mux2_1 _19581_ (.A0(\rbzero.pov.ready_buffer[60] ),
    .A1(_07432_),
    .S(_02963_),
    .X(_02964_));
 sky130_fd_sc_hd__nand2_1 _19582_ (.A(_07431_),
    .B(_02960_),
    .Y(_02965_));
 sky130_fd_sc_hd__o211a_1 _19583_ (.A1(_02956_),
    .A2(_02964_),
    .B1(_02965_),
    .C1(_02780_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _19584_ (.A0(\rbzero.pov.ready_buffer[61] ),
    .A1(_07464_),
    .S(_02963_),
    .X(_02966_));
 sky130_fd_sc_hd__nand2_1 _19585_ (.A(_07462_),
    .B(_02960_),
    .Y(_02967_));
 sky130_fd_sc_hd__o211a_1 _19586_ (.A1(_02956_),
    .A2(_02966_),
    .B1(_02967_),
    .C1(_02780_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _19587_ (.A0(\rbzero.pov.ready_buffer[62] ),
    .A1(_07367_),
    .S(_02963_),
    .X(_02968_));
 sky130_fd_sc_hd__nand2_1 _19588_ (.A(_07340_),
    .B(_02960_),
    .Y(_02969_));
 sky130_fd_sc_hd__o211a_1 _19589_ (.A1(_02956_),
    .A2(_02968_),
    .B1(_02969_),
    .C1(_02780_),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _19590_ (.A0(\rbzero.pov.ready_buffer[63] ),
    .A1(_07395_),
    .S(_02962_),
    .X(_02970_));
 sky130_fd_sc_hd__nand2_1 _19591_ (.A(_07394_),
    .B(_02960_),
    .Y(_02971_));
 sky130_fd_sc_hd__o211a_1 _19592_ (.A1(_02956_),
    .A2(_02970_),
    .B1(_02971_),
    .C1(_02780_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _19593_ (.A0(\rbzero.pov.ready_buffer[64] ),
    .A1(_07413_),
    .S(_02962_),
    .X(_02972_));
 sky130_fd_sc_hd__nand2_1 _19594_ (.A(_07410_),
    .B(_02960_),
    .Y(_02973_));
 sky130_fd_sc_hd__o211a_1 _19595_ (.A1(_02956_),
    .A2(_02972_),
    .B1(_02973_),
    .C1(_02780_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _19596_ (.A0(\rbzero.pov.ready_buffer[65] ),
    .A1(_07539_),
    .S(_02962_),
    .X(_02974_));
 sky130_fd_sc_hd__nand2_1 _19597_ (.A(_07537_),
    .B(_02960_),
    .Y(_02975_));
 sky130_fd_sc_hd__o211a_1 _19598_ (.A1(_02956_),
    .A2(_02974_),
    .B1(_02975_),
    .C1(_02780_),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _19599_ (.A0(\rbzero.pov.ready_buffer[66] ),
    .A1(_07546_),
    .S(_02962_),
    .X(_02976_));
 sky130_fd_sc_hd__nand2_1 _19600_ (.A(_07493_),
    .B(_02960_),
    .Y(_02977_));
 sky130_fd_sc_hd__buf_2 _19601_ (.A(_02727_),
    .X(_02978_));
 sky130_fd_sc_hd__o211a_1 _19602_ (.A1(_02956_),
    .A2(_02976_),
    .B1(_02977_),
    .C1(_02978_),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _19603_ (.A0(\rbzero.pov.ready_buffer[67] ),
    .A1(_07564_),
    .S(_02962_),
    .X(_02979_));
 sky130_fd_sc_hd__nand2_1 _19604_ (.A(_07494_),
    .B(_02955_),
    .Y(_02980_));
 sky130_fd_sc_hd__o211a_1 _19605_ (.A1(_02956_),
    .A2(_02979_),
    .B1(_02980_),
    .C1(_02978_),
    .X(_00968_));
 sky130_fd_sc_hd__o21a_1 _19606_ (.A1(net39),
    .A2(_02954_),
    .B1(_02720_),
    .X(_02981_));
 sky130_fd_sc_hd__or2_1 _19607_ (.A(\rbzero.debug_overlay.playerX[0] ),
    .B(_07562_),
    .X(_02982_));
 sky130_fd_sc_hd__nand2_1 _19608_ (.A(\rbzero.debug_overlay.playerX[0] ),
    .B(_07562_),
    .Y(_02983_));
 sky130_fd_sc_hd__a21oi_1 _19609_ (.A1(_02982_),
    .A2(_02983_),
    .B1(_02835_),
    .Y(_02984_));
 sky130_fd_sc_hd__a211o_1 _19610_ (.A1(\rbzero.pov.ready_buffer[68] ),
    .A2(_02836_),
    .B1(_02955_),
    .C1(_02984_),
    .X(_02985_));
 sky130_fd_sc_hd__o211a_1 _19611_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_02981_),
    .B1(_02985_),
    .C1(_02978_),
    .X(_00969_));
 sky130_fd_sc_hd__o21ai_1 _19612_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_02982_),
    .B1(_02962_),
    .Y(_02986_));
 sky130_fd_sc_hd__a21o_1 _19613_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_02982_),
    .B1(_02986_),
    .X(_02987_));
 sky130_fd_sc_hd__o211a_1 _19614_ (.A1(\rbzero.pov.ready_buffer[69] ),
    .A2(_02963_),
    .B1(_02981_),
    .C1(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__buf_4 _19615_ (.A(_02753_),
    .X(_02989_));
 sky130_fd_sc_hd__a211o_1 _19616_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_02956_),
    .B1(_02988_),
    .C1(_02989_),
    .X(_00970_));
 sky130_fd_sc_hd__o21a_1 _19617_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_02982_),
    .B1(\rbzero.debug_overlay.playerX[2] ),
    .X(_02990_));
 sky130_fd_sc_hd__or3_1 _19618_ (.A(\rbzero.debug_overlay.playerX[2] ),
    .B(\rbzero.debug_overlay.playerX[1] ),
    .C(_02982_),
    .X(_02991_));
 sky130_fd_sc_hd__or3b_1 _19619_ (.A(_02990_),
    .B(_02835_),
    .C_N(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__o211a_1 _19620_ (.A1(\rbzero.pov.ready_buffer[70] ),
    .A2(_02963_),
    .B1(_02981_),
    .C1(_02992_),
    .X(_02993_));
 sky130_fd_sc_hd__a211o_1 _19621_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_02960_),
    .B1(_02993_),
    .C1(_02989_),
    .X(_00971_));
 sky130_fd_sc_hd__and2_1 _19622_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .B(_02991_),
    .X(_02994_));
 sky130_fd_sc_hd__nor2_1 _19623_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .B(_02991_),
    .Y(_02995_));
 sky130_fd_sc_hd__or3_1 _19624_ (.A(_02834_),
    .B(_02994_),
    .C(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__o211a_1 _19625_ (.A1(\rbzero.pov.ready_buffer[71] ),
    .A2(_02963_),
    .B1(_02981_),
    .C1(_02996_),
    .X(_02997_));
 sky130_fd_sc_hd__a211o_1 _19626_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_02960_),
    .B1(_02997_),
    .C1(_02989_),
    .X(_00972_));
 sky130_fd_sc_hd__nor2_1 _19627_ (.A(_02833_),
    .B(_02995_),
    .Y(_02998_));
 sky130_fd_sc_hd__o21ai_1 _19628_ (.A1(_02955_),
    .A2(_02998_),
    .B1(\rbzero.debug_overlay.playerX[4] ),
    .Y(_02999_));
 sky130_fd_sc_hd__and2b_1 _19629_ (.A_N(\rbzero.debug_overlay.playerX[4] ),
    .B(_02995_),
    .X(_03000_));
 sky130_fd_sc_hd__o21a_1 _19630_ (.A1(_02833_),
    .A2(_03000_),
    .B1(_02981_),
    .X(_03001_));
 sky130_fd_sc_hd__o21ai_1 _19631_ (.A1(\rbzero.pov.ready_buffer[72] ),
    .A2(_02963_),
    .B1(_03001_),
    .Y(_03002_));
 sky130_fd_sc_hd__buf_4 _19632_ (.A(_02753_),
    .X(_03003_));
 sky130_fd_sc_hd__a21oi_1 _19633_ (.A1(_02999_),
    .A2(_03002_),
    .B1(_03003_),
    .Y(_00973_));
 sky130_fd_sc_hd__or2_1 _19634_ (.A(\rbzero.debug_overlay.playerX[5] ),
    .B(_03001_),
    .X(_03004_));
 sky130_fd_sc_hd__a21oi_1 _19635_ (.A1(\rbzero.debug_overlay.playerX[5] ),
    .A2(_03000_),
    .B1(_02835_),
    .Y(_03005_));
 sky130_fd_sc_hd__a211o_1 _19636_ (.A1(\rbzero.pov.ready_buffer[73] ),
    .A2(_02836_),
    .B1(_02955_),
    .C1(_03005_),
    .X(_03006_));
 sky130_fd_sc_hd__a21o_1 _19637_ (.A1(_03004_),
    .A2(_03006_),
    .B1(_03003_),
    .X(_00974_));
 sky130_fd_sc_hd__o21ai_2 _19638_ (.A1(net40),
    .A2(_02954_),
    .B1(_02721_),
    .Y(_03007_));
 sky130_fd_sc_hd__buf_2 _19639_ (.A(_03007_),
    .X(_03008_));
 sky130_fd_sc_hd__inv_2 _19640_ (.A(\rbzero.debug_overlay.playerY[-9] ),
    .Y(_03009_));
 sky130_fd_sc_hd__mux2_1 _19641_ (.A0(_03009_),
    .A1(\rbzero.pov.ready_buffer[44] ),
    .S(_02835_),
    .X(_03010_));
 sky130_fd_sc_hd__nand2_1 _19642_ (.A(_03009_),
    .B(_03008_),
    .Y(_03011_));
 sky130_fd_sc_hd__o211a_1 _19643_ (.A1(_03008_),
    .A2(_03010_),
    .B1(_03011_),
    .C1(_02978_),
    .X(_00975_));
 sky130_fd_sc_hd__o21a_2 _19644_ (.A1(net40),
    .A2(_02954_),
    .B1(_02721_),
    .X(_03012_));
 sky130_fd_sc_hd__nand2_1 _19645_ (.A(\rbzero.pov.ready_buffer[45] ),
    .B(_02835_),
    .Y(_03013_));
 sky130_fd_sc_hd__o211a_1 _19646_ (.A1(_07427_),
    .A2(_02835_),
    .B1(_03012_),
    .C1(_03013_),
    .X(_03014_));
 sky130_fd_sc_hd__buf_4 _19647_ (.A(_03442_),
    .X(_03015_));
 sky130_fd_sc_hd__a211oi_1 _19648_ (.A1(_08574_),
    .A2(_03008_),
    .B1(_03014_),
    .C1(_03015_),
    .Y(_00976_));
 sky130_fd_sc_hd__buf_2 _19649_ (.A(_03012_),
    .X(_03016_));
 sky130_fd_sc_hd__nor2_1 _19650_ (.A(_07458_),
    .B(_02958_),
    .Y(_03017_));
 sky130_fd_sc_hd__a211o_1 _19651_ (.A1(\rbzero.pov.ready_buffer[46] ),
    .A2(_02836_),
    .B1(_03008_),
    .C1(_03017_),
    .X(_03018_));
 sky130_fd_sc_hd__o211a_1 _19652_ (.A1(\rbzero.debug_overlay.playerY[-7] ),
    .A2(_03016_),
    .B1(_03018_),
    .C1(_02978_),
    .X(_00977_));
 sky130_fd_sc_hd__nor2_1 _19653_ (.A(_07360_),
    .B(_02958_),
    .Y(_03019_));
 sky130_fd_sc_hd__a211o_1 _19654_ (.A1(\rbzero.pov.ready_buffer[47] ),
    .A2(_02836_),
    .B1(_03008_),
    .C1(_03019_),
    .X(_03020_));
 sky130_fd_sc_hd__o211a_1 _19655_ (.A1(\rbzero.debug_overlay.playerY[-6] ),
    .A2(_03016_),
    .B1(_03020_),
    .C1(_02978_),
    .X(_00978_));
 sky130_fd_sc_hd__nor2_1 _19656_ (.A(_07390_),
    .B(_02958_),
    .Y(_03021_));
 sky130_fd_sc_hd__a211o_1 _19657_ (.A1(\rbzero.pov.ready_buffer[48] ),
    .A2(_02836_),
    .B1(_03008_),
    .C1(_03021_),
    .X(_03022_));
 sky130_fd_sc_hd__o211a_1 _19658_ (.A1(\rbzero.debug_overlay.playerY[-5] ),
    .A2(_03016_),
    .B1(_03022_),
    .C1(_02978_),
    .X(_00979_));
 sky130_fd_sc_hd__nor2_1 _19659_ (.A(_07406_),
    .B(_02958_),
    .Y(_03023_));
 sky130_fd_sc_hd__a211o_1 _19660_ (.A1(\rbzero.pov.ready_buffer[49] ),
    .A2(_02958_),
    .B1(_03008_),
    .C1(_03023_),
    .X(_03024_));
 sky130_fd_sc_hd__o211a_1 _19661_ (.A1(\rbzero.debug_overlay.playerY[-4] ),
    .A2(_03016_),
    .B1(_03024_),
    .C1(_02978_),
    .X(_00980_));
 sky130_fd_sc_hd__nor2_1 _19662_ (.A(_07534_),
    .B(_02958_),
    .Y(_03025_));
 sky130_fd_sc_hd__a211o_1 _19663_ (.A1(\rbzero.pov.ready_buffer[50] ),
    .A2(_02958_),
    .B1(_03007_),
    .C1(_03025_),
    .X(_03026_));
 sky130_fd_sc_hd__o211a_1 _19664_ (.A1(\rbzero.debug_overlay.playerY[-3] ),
    .A2(_03016_),
    .B1(_03026_),
    .C1(_02978_),
    .X(_00981_));
 sky130_fd_sc_hd__nand2_1 _19665_ (.A(\rbzero.pov.ready_buffer[51] ),
    .B(_02836_),
    .Y(_03027_));
 sky130_fd_sc_hd__o211ai_1 _19666_ (.A1(_07543_),
    .A2(_02836_),
    .B1(_03016_),
    .C1(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__o211a_1 _19667_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_03016_),
    .B1(_03028_),
    .C1(_02978_),
    .X(_00982_));
 sky130_fd_sc_hd__nand2_1 _19668_ (.A(\rbzero.pov.ready_buffer[52] ),
    .B(_02836_),
    .Y(_03029_));
 sky130_fd_sc_hd__o211ai_1 _19669_ (.A1(_07558_),
    .A2(_02836_),
    .B1(_03012_),
    .C1(_03029_),
    .Y(_03030_));
 sky130_fd_sc_hd__buf_4 _19670_ (.A(_02727_),
    .X(_03031_));
 sky130_fd_sc_hd__o211a_1 _19671_ (.A1(\rbzero.debug_overlay.playerY[-1] ),
    .A2(_03016_),
    .B1(_03030_),
    .C1(_03031_),
    .X(_00983_));
 sky130_fd_sc_hd__or2_1 _19672_ (.A(\rbzero.debug_overlay.playerY[0] ),
    .B(_07498_),
    .X(_03032_));
 sky130_fd_sc_hd__nand2_1 _19673_ (.A(\rbzero.debug_overlay.playerY[0] ),
    .B(_07498_),
    .Y(_03033_));
 sky130_fd_sc_hd__a21oi_1 _19674_ (.A1(_03032_),
    .A2(_03033_),
    .B1(_02835_),
    .Y(_03034_));
 sky130_fd_sc_hd__a211o_1 _19675_ (.A1(\rbzero.pov.ready_buffer[53] ),
    .A2(_02958_),
    .B1(_03007_),
    .C1(_03034_),
    .X(_03035_));
 sky130_fd_sc_hd__o211a_1 _19676_ (.A1(\rbzero.debug_overlay.playerY[0] ),
    .A2(_03016_),
    .B1(_03035_),
    .C1(_03031_),
    .X(_00984_));
 sky130_fd_sc_hd__o21ai_1 _19677_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_03032_),
    .B1(_02962_),
    .Y(_03036_));
 sky130_fd_sc_hd__a21o_1 _19678_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_03032_),
    .B1(_03036_),
    .X(_03037_));
 sky130_fd_sc_hd__o211a_1 _19679_ (.A1(\rbzero.pov.ready_buffer[54] ),
    .A2(_02963_),
    .B1(_03012_),
    .C1(_03037_),
    .X(_03038_));
 sky130_fd_sc_hd__a211o_1 _19680_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_03008_),
    .B1(_03038_),
    .C1(_02989_),
    .X(_00985_));
 sky130_fd_sc_hd__or3_1 _19681_ (.A(\rbzero.debug_overlay.playerY[2] ),
    .B(\rbzero.debug_overlay.playerY[1] ),
    .C(_03032_),
    .X(_03039_));
 sky130_fd_sc_hd__o21ai_1 _19682_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_03032_),
    .B1(\rbzero.debug_overlay.playerY[2] ),
    .Y(_03040_));
 sky130_fd_sc_hd__a21oi_1 _19683_ (.A1(_03039_),
    .A2(_03040_),
    .B1(_02835_),
    .Y(_03041_));
 sky130_fd_sc_hd__a211o_1 _19684_ (.A1(\rbzero.pov.ready_buffer[55] ),
    .A2(_02958_),
    .B1(_03007_),
    .C1(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__o211a_1 _19685_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_03016_),
    .B1(_03042_),
    .C1(_03031_),
    .X(_00986_));
 sky130_fd_sc_hd__or2_1 _19686_ (.A(\rbzero.debug_overlay.playerY[3] ),
    .B(_03039_),
    .X(_03043_));
 sky130_fd_sc_hd__inv_2 _19687_ (.A(_03043_),
    .Y(_03044_));
 sky130_fd_sc_hd__a21o_1 _19688_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_03039_),
    .B1(_02835_),
    .X(_03045_));
 sky130_fd_sc_hd__o221a_1 _19689_ (.A1(\rbzero.pov.ready_buffer[56] ),
    .A2(_02963_),
    .B1(_03044_),
    .B2(_03045_),
    .C1(_03012_),
    .X(_03046_));
 sky130_fd_sc_hd__a211o_1 _19690_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_03008_),
    .B1(_03046_),
    .C1(_02989_),
    .X(_00987_));
 sky130_fd_sc_hd__nor2_1 _19691_ (.A(_02833_),
    .B(_03044_),
    .Y(_03047_));
 sky130_fd_sc_hd__o21ai_1 _19692_ (.A1(_03008_),
    .A2(_03047_),
    .B1(\rbzero.debug_overlay.playerY[4] ),
    .Y(_03048_));
 sky130_fd_sc_hd__nor2_1 _19693_ (.A(\rbzero.debug_overlay.playerY[4] ),
    .B(_03043_),
    .Y(_03049_));
 sky130_fd_sc_hd__o21a_1 _19694_ (.A1(_02833_),
    .A2(_03049_),
    .B1(_03012_),
    .X(_03050_));
 sky130_fd_sc_hd__o21ai_1 _19695_ (.A1(\rbzero.pov.ready_buffer[57] ),
    .A2(_02963_),
    .B1(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__a21oi_1 _19696_ (.A1(_03048_),
    .A2(_03051_),
    .B1(_03003_),
    .Y(_00988_));
 sky130_fd_sc_hd__or4b_1 _19697_ (.A(\rbzero.debug_overlay.playerY[4] ),
    .B(_02834_),
    .C(_03043_),
    .D_N(\rbzero.debug_overlay.playerY[5] ),
    .X(_03052_));
 sky130_fd_sc_hd__o21ai_1 _19698_ (.A1(\rbzero.pov.ready_buffer[58] ),
    .A2(_02962_),
    .B1(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__a2bb2o_1 _19699_ (.A1_N(\rbzero.debug_overlay.playerY[5] ),
    .A2_N(_03050_),
    .B1(_03053_),
    .B2(_03012_),
    .X(_03054_));
 sky130_fd_sc_hd__nand2_1 _19700_ (.A(_02728_),
    .B(_03054_),
    .Y(_00989_));
 sky130_fd_sc_hd__nand3_2 _19701_ (.A(\rbzero.pov.ready ),
    .B(_02721_),
    .C(_02833_),
    .Y(_03055_));
 sky130_fd_sc_hd__buf_2 _19702_ (.A(_03055_),
    .X(_03056_));
 sky130_fd_sc_hd__and3_1 _19703_ (.A(\rbzero.pov.ready ),
    .B(_02720_),
    .C(_02833_),
    .X(_03057_));
 sky130_fd_sc_hd__clkbuf_2 _19704_ (.A(_03057_),
    .X(_03058_));
 sky130_fd_sc_hd__buf_2 _19705_ (.A(_03058_),
    .X(_03059_));
 sky130_fd_sc_hd__o221a_1 _19706_ (.A1(\rbzero.pov.ready_buffer[33] ),
    .A2(_03056_),
    .B1(_03059_),
    .B2(\rbzero.debug_overlay.facingX[-9] ),
    .C1(_03031_),
    .X(_00990_));
 sky130_fd_sc_hd__and3_1 _19707_ (.A(\rbzero.pov.ready ),
    .B(_02721_),
    .C(_02833_),
    .X(_03060_));
 sky130_fd_sc_hd__buf_2 _19708_ (.A(_03060_),
    .X(_03061_));
 sky130_fd_sc_hd__nand2_1 _19709_ (.A(_02721_),
    .B(_02954_),
    .Y(_03062_));
 sky130_fd_sc_hd__buf_2 _19710_ (.A(_03062_),
    .X(_03063_));
 sky130_fd_sc_hd__buf_4 _19711_ (.A(_02708_),
    .X(_03064_));
 sky130_fd_sc_hd__a221o_1 _19712_ (.A1(\rbzero.pov.ready_buffer[34] ),
    .A2(_03061_),
    .B1(_03063_),
    .B2(\rbzero.debug_overlay.facingX[-8] ),
    .C1(_03064_),
    .X(_00991_));
 sky130_fd_sc_hd__o221a_1 _19713_ (.A1(\rbzero.pov.ready_buffer[35] ),
    .A2(_03056_),
    .B1(_03059_),
    .B2(\rbzero.debug_overlay.facingX[-7] ),
    .C1(_03031_),
    .X(_00992_));
 sky130_fd_sc_hd__o221a_1 _19714_ (.A1(\rbzero.pov.ready_buffer[36] ),
    .A2(_03056_),
    .B1(_03059_),
    .B2(\rbzero.debug_overlay.facingX[-6] ),
    .C1(_03031_),
    .X(_00993_));
 sky130_fd_sc_hd__o221a_1 _19715_ (.A1(\rbzero.pov.ready_buffer[37] ),
    .A2(_03056_),
    .B1(_03059_),
    .B2(\rbzero.debug_overlay.facingX[-5] ),
    .C1(_03031_),
    .X(_00994_));
 sky130_fd_sc_hd__buf_2 _19716_ (.A(_02727_),
    .X(_03065_));
 sky130_fd_sc_hd__o221a_1 _19717_ (.A1(\rbzero.pov.ready_buffer[38] ),
    .A2(_03056_),
    .B1(_03059_),
    .B2(\rbzero.debug_overlay.facingX[-4] ),
    .C1(_03065_),
    .X(_00995_));
 sky130_fd_sc_hd__a221o_1 _19718_ (.A1(\rbzero.pov.ready_buffer[39] ),
    .A2(_03061_),
    .B1(_03063_),
    .B2(\rbzero.debug_overlay.facingX[-3] ),
    .C1(_03064_),
    .X(_00996_));
 sky130_fd_sc_hd__buf_2 _19719_ (.A(_02708_),
    .X(_03066_));
 sky130_fd_sc_hd__a221o_1 _19720_ (.A1(\rbzero.pov.ready_buffer[40] ),
    .A2(_03061_),
    .B1(_03063_),
    .B2(\rbzero.debug_overlay.facingX[-2] ),
    .C1(_03066_),
    .X(_00997_));
 sky130_fd_sc_hd__a221o_1 _19721_ (.A1(\rbzero.pov.ready_buffer[41] ),
    .A2(_03061_),
    .B1(_03063_),
    .B2(\rbzero.debug_overlay.facingX[-1] ),
    .C1(_03066_),
    .X(_00998_));
 sky130_fd_sc_hd__o221a_1 _19722_ (.A1(\rbzero.pov.ready_buffer[42] ),
    .A2(_03056_),
    .B1(_03059_),
    .B2(\rbzero.debug_overlay.facingX[0] ),
    .C1(_03065_),
    .X(_00999_));
 sky130_fd_sc_hd__a221o_1 _19723_ (.A1(\rbzero.pov.ready_buffer[43] ),
    .A2(_03061_),
    .B1(_03063_),
    .B2(\rbzero.debug_overlay.facingX[10] ),
    .C1(_03066_),
    .X(_01000_));
 sky130_fd_sc_hd__a221o_1 _19724_ (.A1(\rbzero.pov.ready_buffer[22] ),
    .A2(_03061_),
    .B1(_03063_),
    .B2(\rbzero.debug_overlay.facingY[-9] ),
    .C1(_03066_),
    .X(_01001_));
 sky130_fd_sc_hd__a221o_1 _19725_ (.A1(\rbzero.pov.ready_buffer[23] ),
    .A2(_03061_),
    .B1(_03063_),
    .B2(\rbzero.debug_overlay.facingY[-8] ),
    .C1(_03066_),
    .X(_01002_));
 sky130_fd_sc_hd__o221a_1 _19726_ (.A1(\rbzero.pov.ready_buffer[24] ),
    .A2(_03056_),
    .B1(_03059_),
    .B2(\rbzero.debug_overlay.facingY[-7] ),
    .C1(_03065_),
    .X(_01003_));
 sky130_fd_sc_hd__o221a_1 _19727_ (.A1(\rbzero.pov.ready_buffer[25] ),
    .A2(_03056_),
    .B1(_03059_),
    .B2(\rbzero.debug_overlay.facingY[-6] ),
    .C1(_03065_),
    .X(_01004_));
 sky130_fd_sc_hd__a221o_1 _19728_ (.A1(\rbzero.pov.ready_buffer[26] ),
    .A2(_03061_),
    .B1(_03063_),
    .B2(\rbzero.debug_overlay.facingY[-5] ),
    .C1(_03066_),
    .X(_01005_));
 sky130_fd_sc_hd__a221o_1 _19729_ (.A1(\rbzero.pov.ready_buffer[27] ),
    .A2(_03061_),
    .B1(_03063_),
    .B2(\rbzero.debug_overlay.facingY[-4] ),
    .C1(_03066_),
    .X(_01006_));
 sky130_fd_sc_hd__a221o_1 _19730_ (.A1(\rbzero.pov.ready_buffer[28] ),
    .A2(_03061_),
    .B1(_03063_),
    .B2(\rbzero.debug_overlay.facingY[-3] ),
    .C1(_03066_),
    .X(_01007_));
 sky130_fd_sc_hd__o221a_1 _19731_ (.A1(\rbzero.pov.ready_buffer[29] ),
    .A2(_03056_),
    .B1(_03059_),
    .B2(\rbzero.debug_overlay.facingY[-2] ),
    .C1(_03065_),
    .X(_01008_));
 sky130_fd_sc_hd__o221a_1 _19732_ (.A1(\rbzero.pov.ready_buffer[30] ),
    .A2(_03056_),
    .B1(_03059_),
    .B2(\rbzero.debug_overlay.facingY[-1] ),
    .C1(_03065_),
    .X(_01009_));
 sky130_fd_sc_hd__buf_2 _19733_ (.A(_03060_),
    .X(_03067_));
 sky130_fd_sc_hd__buf_2 _19734_ (.A(_03062_),
    .X(_03068_));
 sky130_fd_sc_hd__a221o_1 _19735_ (.A1(\rbzero.pov.ready_buffer[31] ),
    .A2(_03067_),
    .B1(_03068_),
    .B2(\rbzero.debug_overlay.facingY[0] ),
    .C1(_03066_),
    .X(_01010_));
 sky130_fd_sc_hd__clkbuf_4 _19736_ (.A(_03055_),
    .X(_03069_));
 sky130_fd_sc_hd__clkbuf_4 _19737_ (.A(_03058_),
    .X(_03070_));
 sky130_fd_sc_hd__o221a_1 _19738_ (.A1(\rbzero.pov.ready_buffer[32] ),
    .A2(_03069_),
    .B1(_03070_),
    .B2(\rbzero.debug_overlay.facingY[10] ),
    .C1(_03065_),
    .X(_01011_));
 sky130_fd_sc_hd__o221a_1 _19739_ (.A1(\rbzero.pov.ready_buffer[11] ),
    .A2(_03069_),
    .B1(_03070_),
    .B2(\rbzero.debug_overlay.vplaneX[-9] ),
    .C1(_03065_),
    .X(_01012_));
 sky130_fd_sc_hd__a221o_1 _19740_ (.A1(\rbzero.pov.ready_buffer[12] ),
    .A2(_03067_),
    .B1(_03068_),
    .B2(\rbzero.debug_overlay.vplaneX[-8] ),
    .C1(_03066_),
    .X(_01013_));
 sky130_fd_sc_hd__a221o_1 _19741_ (.A1(\rbzero.pov.ready_buffer[13] ),
    .A2(_03067_),
    .B1(_03068_),
    .B2(\rbzero.debug_overlay.vplaneX[-7] ),
    .C1(_03015_),
    .X(_01014_));
 sky130_fd_sc_hd__o221a_1 _19742_ (.A1(\rbzero.pov.ready_buffer[14] ),
    .A2(_03069_),
    .B1(_03070_),
    .B2(\rbzero.debug_overlay.vplaneX[-6] ),
    .C1(_03065_),
    .X(_01015_));
 sky130_fd_sc_hd__o221a_1 _19743_ (.A1(\rbzero.pov.ready_buffer[15] ),
    .A2(_03069_),
    .B1(_03070_),
    .B2(\rbzero.debug_overlay.vplaneX[-5] ),
    .C1(_03065_),
    .X(_01016_));
 sky130_fd_sc_hd__o221a_1 _19744_ (.A1(\rbzero.pov.ready_buffer[16] ),
    .A2(_03069_),
    .B1(_03070_),
    .B2(\rbzero.debug_overlay.vplaneX[-4] ),
    .C1(_02832_),
    .X(_01017_));
 sky130_fd_sc_hd__a221o_1 _19745_ (.A1(\rbzero.pov.ready_buffer[17] ),
    .A2(_03067_),
    .B1(_03068_),
    .B2(\rbzero.debug_overlay.vplaneX[-3] ),
    .C1(_03015_),
    .X(_01018_));
 sky130_fd_sc_hd__a221o_1 _19746_ (.A1(\rbzero.pov.ready_buffer[18] ),
    .A2(_03067_),
    .B1(_03068_),
    .B2(\rbzero.debug_overlay.vplaneX[-2] ),
    .C1(_03015_),
    .X(_01019_));
 sky130_fd_sc_hd__o221a_1 _19747_ (.A1(\rbzero.pov.ready_buffer[19] ),
    .A2(_03069_),
    .B1(_03070_),
    .B2(_02191_),
    .C1(_02832_),
    .X(_01020_));
 sky130_fd_sc_hd__a221o_1 _19748_ (.A1(\rbzero.pov.ready_buffer[20] ),
    .A2(_03067_),
    .B1(_03068_),
    .B2(\rbzero.debug_overlay.vplaneX[0] ),
    .C1(_03015_),
    .X(_01021_));
 sky130_fd_sc_hd__o221a_1 _19749_ (.A1(\rbzero.pov.ready_buffer[21] ),
    .A2(_03069_),
    .B1(_03070_),
    .B2(_02275_),
    .C1(_02832_),
    .X(_01022_));
 sky130_fd_sc_hd__a221o_1 _19750_ (.A1(\rbzero.pov.ready_buffer[0] ),
    .A2(_03067_),
    .B1(_03068_),
    .B2(\rbzero.debug_overlay.vplaneY[-9] ),
    .C1(_03015_),
    .X(_01023_));
 sky130_fd_sc_hd__o221a_1 _19751_ (.A1(\rbzero.pov.ready_buffer[1] ),
    .A2(_03069_),
    .B1(_03070_),
    .B2(\rbzero.debug_overlay.vplaneY[-8] ),
    .C1(_02832_),
    .X(_01024_));
 sky130_fd_sc_hd__o221a_1 _19752_ (.A1(\rbzero.pov.ready_buffer[2] ),
    .A2(_03069_),
    .B1(_03070_),
    .B2(\rbzero.debug_overlay.vplaneY[-7] ),
    .C1(_02832_),
    .X(_01025_));
 sky130_fd_sc_hd__o221a_1 _19753_ (.A1(\rbzero.pov.ready_buffer[3] ),
    .A2(_03069_),
    .B1(_03070_),
    .B2(\rbzero.debug_overlay.vplaneY[-6] ),
    .C1(_02832_),
    .X(_01026_));
 sky130_fd_sc_hd__o221a_1 _19754_ (.A1(\rbzero.pov.ready_buffer[4] ),
    .A2(_03055_),
    .B1(_03058_),
    .B2(\rbzero.debug_overlay.vplaneY[-5] ),
    .C1(_02832_),
    .X(_01027_));
 sky130_fd_sc_hd__a221o_1 _19755_ (.A1(\rbzero.pov.ready_buffer[5] ),
    .A2(_03067_),
    .B1(_03068_),
    .B2(\rbzero.debug_overlay.vplaneY[-4] ),
    .C1(_03015_),
    .X(_01028_));
 sky130_fd_sc_hd__a221o_1 _19756_ (.A1(\rbzero.pov.ready_buffer[6] ),
    .A2(_03067_),
    .B1(_03068_),
    .B2(\rbzero.debug_overlay.vplaneY[-3] ),
    .C1(_03015_),
    .X(_01029_));
 sky130_fd_sc_hd__a221o_1 _19757_ (.A1(\rbzero.pov.ready_buffer[7] ),
    .A2(_03067_),
    .B1(_03068_),
    .B2(_04260_),
    .C1(_03015_),
    .X(_01030_));
 sky130_fd_sc_hd__o221a_1 _19758_ (.A1(\rbzero.pov.ready_buffer[8] ),
    .A2(_03055_),
    .B1(_03058_),
    .B2(\rbzero.debug_overlay.vplaneY[-1] ),
    .C1(_02832_),
    .X(_01031_));
 sky130_fd_sc_hd__a221o_1 _19759_ (.A1(\rbzero.pov.ready_buffer[9] ),
    .A2(_03060_),
    .B1(_03062_),
    .B2(_02428_),
    .C1(_03015_),
    .X(_01032_));
 sky130_fd_sc_hd__o221a_1 _19760_ (.A1(\rbzero.pov.ready_buffer[10] ),
    .A2(_03055_),
    .B1(_03058_),
    .B2(_02510_),
    .C1(_02832_),
    .X(_01033_));
 sky130_fd_sc_hd__a31o_1 _19761_ (.A1(_02838_),
    .A2(_02837_),
    .A3(_02843_),
    .B1(\rbzero.pov.spi_done ),
    .X(_03071_));
 sky130_fd_sc_hd__and2_1 _19762_ (.A(_02608_),
    .B(_03071_),
    .X(_03072_));
 sky130_fd_sc_hd__clkbuf_1 _19763_ (.A(_03072_),
    .X(_01034_));
 sky130_fd_sc_hd__inv_2 _19764_ (.A(_04632_),
    .Y(_03073_));
 sky130_fd_sc_hd__or4_1 _19765_ (.A(_04110_),
    .B(_04106_),
    .C(_03073_),
    .D(_04114_),
    .X(_03074_));
 sky130_fd_sc_hd__or4_1 _19766_ (.A(_04246_),
    .B(_04628_),
    .C(_04631_),
    .D(_03074_),
    .X(_03075_));
 sky130_fd_sc_hd__or4b_1 _19767_ (.A(_04246_),
    .B(_04632_),
    .C(\gpout0.vpos[0] ),
    .D_N(_04628_),
    .X(_03076_));
 sky130_fd_sc_hd__o41a_1 _19768_ (.A1(_04110_),
    .A2(_04106_),
    .A3(_04114_),
    .A4(_03076_),
    .B1(_04920_),
    .X(_03077_));
 sky130_fd_sc_hd__a21boi_1 _19769_ (.A1(o_vsync),
    .A2(_03075_),
    .B1_N(_03077_),
    .Y(_01035_));
 sky130_fd_sc_hd__or4b_1 _19770_ (.A(_04080_),
    .B(_04591_),
    .C(_04592_),
    .D_N(_04078_),
    .X(_03078_));
 sky130_fd_sc_hd__or4_1 _19771_ (.A(_03289_),
    .B(_03443_),
    .C(_03803_),
    .D(_03078_),
    .X(_03079_));
 sky130_fd_sc_hd__nand2_1 _19772_ (.A(_03784_),
    .B(_03781_),
    .Y(_03080_));
 sky130_fd_sc_hd__o41a_1 _19773_ (.A1(_03289_),
    .A2(_03443_),
    .A3(_03080_),
    .A4(_03078_),
    .B1(_04920_),
    .X(_03081_));
 sky130_fd_sc_hd__a21boi_1 _19774_ (.A1(o_hsync),
    .A2(_03079_),
    .B1_N(_03081_),
    .Y(_01036_));
 sky130_fd_sc_hd__or4_1 _19775_ (.A(_04111_),
    .B(\gpout0.vpos[6] ),
    .C(_04104_),
    .D(_04106_),
    .X(_03082_));
 sky130_fd_sc_hd__or4_1 _19776_ (.A(\gpout0.vpos[8] ),
    .B(\gpout0.vpos[7] ),
    .C(_03076_),
    .D(_03082_),
    .X(_03083_));
 sky130_fd_sc_hd__inv_2 _19777_ (.A(_03083_),
    .Y(_03084_));
 sky130_fd_sc_hd__nor2_1 _19778_ (.A(_03813_),
    .B(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__nand2_1 _19779_ (.A(_04631_),
    .B(_03808_),
    .Y(_03086_));
 sky130_fd_sc_hd__o211a_1 _19780_ (.A1(_04631_),
    .A2(_03085_),
    .B1(_03086_),
    .C1(_03031_),
    .X(_01037_));
 sky130_fd_sc_hd__a31o_1 _19781_ (.A1(_04632_),
    .A2(_04631_),
    .A3(_03808_),
    .B1(_02753_),
    .X(_03087_));
 sky130_fd_sc_hd__a21oi_1 _19782_ (.A1(_03073_),
    .A2(_03086_),
    .B1(_03087_),
    .Y(_01038_));
 sky130_fd_sc_hd__a22o_1 _19783_ (.A1(_04628_),
    .A2(_03813_),
    .B1(_02717_),
    .B2(_03085_),
    .X(_03088_));
 sky130_fd_sc_hd__a21o_1 _19784_ (.A1(_04632_),
    .A2(_04631_),
    .B1(_04628_),
    .X(_03089_));
 sky130_fd_sc_hd__and3_1 _19785_ (.A(_09247_),
    .B(_03088_),
    .C(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__clkbuf_1 _19786_ (.A(_03090_),
    .X(_01039_));
 sky130_fd_sc_hd__or2_1 _19787_ (.A(_04101_),
    .B(_02716_),
    .X(_03091_));
 sky130_fd_sc_hd__nor2_1 _19788_ (.A(_02753_),
    .B(_02718_),
    .Y(_03092_));
 sky130_fd_sc_hd__clkbuf_4 _19789_ (.A(_09245_),
    .X(_03093_));
 sky130_fd_sc_hd__a32o_1 _19790_ (.A1(_03085_),
    .A2(_03091_),
    .A3(_03092_),
    .B1(_03093_),
    .B2(_04101_),
    .X(_01040_));
 sky130_fd_sc_hd__and3_1 _19791_ (.A(_04106_),
    .B(_03808_),
    .C(_02718_),
    .X(_03094_));
 sky130_fd_sc_hd__o21ai_1 _19792_ (.A1(_04106_),
    .A2(_02719_),
    .B1(_02742_),
    .Y(_03095_));
 sky130_fd_sc_hd__nor2_1 _19793_ (.A(_03094_),
    .B(_03095_),
    .Y(_01041_));
 sky130_fd_sc_hd__and2_1 _19794_ (.A(_04104_),
    .B(_03094_),
    .X(_03096_));
 sky130_fd_sc_hd__o21ai_1 _19795_ (.A1(_04104_),
    .A2(_03094_),
    .B1(_02742_),
    .Y(_03097_));
 sky130_fd_sc_hd__nor2_1 _19796_ (.A(_03096_),
    .B(_03097_),
    .Y(_01042_));
 sky130_fd_sc_hd__nand2_1 _19797_ (.A(\gpout0.vpos[6] ),
    .B(_03096_),
    .Y(_03098_));
 sky130_fd_sc_hd__o211a_1 _19798_ (.A1(\gpout0.vpos[6] ),
    .A2(_03096_),
    .B1(_03098_),
    .C1(_03031_),
    .X(_01043_));
 sky130_fd_sc_hd__and3_1 _19799_ (.A(\gpout0.vpos[7] ),
    .B(\gpout0.vpos[6] ),
    .C(_03096_),
    .X(_03099_));
 sky130_fd_sc_hd__a31o_1 _19800_ (.A1(\gpout0.vpos[6] ),
    .A2(_04104_),
    .A3(_03094_),
    .B1(\gpout0.vpos[7] ),
    .X(_03100_));
 sky130_fd_sc_hd__and3b_1 _19801_ (.A_N(_03099_),
    .B(_04920_),
    .C(_03100_),
    .X(_03101_));
 sky130_fd_sc_hd__clkbuf_1 _19802_ (.A(_03101_),
    .X(_01044_));
 sky130_fd_sc_hd__nand2_1 _19803_ (.A(_04113_),
    .B(_03096_),
    .Y(_03102_));
 sky130_fd_sc_hd__o211a_1 _19804_ (.A1(\gpout0.vpos[8] ),
    .A2(_03099_),
    .B1(_03102_),
    .C1(_03031_),
    .X(_01045_));
 sky130_fd_sc_hd__a41o_1 _19805_ (.A1(_04104_),
    .A2(_04106_),
    .A3(_04113_),
    .A4(_02718_),
    .B1(_03084_),
    .X(_03103_));
 sky130_fd_sc_hd__a31o_1 _19806_ (.A1(_04110_),
    .A2(_03808_),
    .A3(_03103_),
    .B1(_02708_),
    .X(_03104_));
 sky130_fd_sc_hd__a21oi_1 _19807_ (.A1(_04111_),
    .A2(_03102_),
    .B1(_03104_),
    .Y(_01046_));
 sky130_fd_sc_hd__a31o_1 _19808_ (.A1(\rbzero.spi_registers.got_new_vinf ),
    .A2(_02742_),
    .A3(_02740_),
    .B1(_02141_),
    .X(_01047_));
 sky130_fd_sc_hd__clkinv_2 _19809_ (.A(_02863_),
    .Y(_00081_));
 sky130_fd_sc_hd__clkinv_2 _19810_ (.A(_02863_),
    .Y(_00082_));
 sky130_fd_sc_hd__clkinv_2 _19811_ (.A(_02863_),
    .Y(_00083_));
 sky130_fd_sc_hd__clkinv_2 _19812_ (.A(_02863_),
    .Y(_00084_));
 sky130_fd_sc_hd__clkinv_2 _19813_ (.A(_02863_),
    .Y(_00085_));
 sky130_fd_sc_hd__clkinv_2 _19814_ (.A(_02863_),
    .Y(_00086_));
 sky130_fd_sc_hd__buf_4 _19815_ (.A(_02862_),
    .X(_03105_));
 sky130_fd_sc_hd__clkinv_2 _19816_ (.A(_03105_),
    .Y(_00087_));
 sky130_fd_sc_hd__clkinv_2 _19817_ (.A(_03105_),
    .Y(_00088_));
 sky130_fd_sc_hd__clkinv_2 _19818_ (.A(_03105_),
    .Y(_00089_));
 sky130_fd_sc_hd__clkinv_2 _19819_ (.A(_03105_),
    .Y(_00090_));
 sky130_fd_sc_hd__clkinv_2 _19820_ (.A(_03105_),
    .Y(_00091_));
 sky130_fd_sc_hd__clkinv_2 _19821_ (.A(_03105_),
    .Y(_00092_));
 sky130_fd_sc_hd__clkinv_2 _19822_ (.A(_03105_),
    .Y(_00093_));
 sky130_fd_sc_hd__clkinv_2 _19823_ (.A(_03105_),
    .Y(_00094_));
 sky130_fd_sc_hd__clkinv_2 _19824_ (.A(_03105_),
    .Y(_00095_));
 sky130_fd_sc_hd__clkinv_2 _19825_ (.A(_03105_),
    .Y(_00096_));
 sky130_fd_sc_hd__buf_4 _19826_ (.A(_02862_),
    .X(_03106_));
 sky130_fd_sc_hd__clkinv_2 _19827_ (.A(_03106_),
    .Y(_00097_));
 sky130_fd_sc_hd__clkinv_2 _19828_ (.A(_03106_),
    .Y(_00098_));
 sky130_fd_sc_hd__clkinv_2 _19829_ (.A(_03106_),
    .Y(_00099_));
 sky130_fd_sc_hd__clkinv_2 _19830_ (.A(_03106_),
    .Y(_00100_));
 sky130_fd_sc_hd__clkinv_2 _19831_ (.A(_03106_),
    .Y(_00101_));
 sky130_fd_sc_hd__clkinv_2 _19832_ (.A(_03106_),
    .Y(_00102_));
 sky130_fd_sc_hd__clkinv_2 _19833_ (.A(_03106_),
    .Y(_00103_));
 sky130_fd_sc_hd__clkinv_2 _19834_ (.A(_03106_),
    .Y(_00104_));
 sky130_fd_sc_hd__clkinv_2 _19835_ (.A(_03106_),
    .Y(_00105_));
 sky130_fd_sc_hd__clkinv_2 _19836_ (.A(_03106_),
    .Y(_00106_));
 sky130_fd_sc_hd__buf_4 _19837_ (.A(_02862_),
    .X(_03107_));
 sky130_fd_sc_hd__clkinv_2 _19838_ (.A(_03107_),
    .Y(_00107_));
 sky130_fd_sc_hd__clkinv_2 _19839_ (.A(_03107_),
    .Y(_00108_));
 sky130_fd_sc_hd__clkinv_2 _19840_ (.A(_03107_),
    .Y(_00109_));
 sky130_fd_sc_hd__clkinv_2 _19841_ (.A(_03107_),
    .Y(_00110_));
 sky130_fd_sc_hd__clkinv_2 _19842_ (.A(_03107_),
    .Y(_00111_));
 sky130_fd_sc_hd__clkinv_2 _19843_ (.A(_03107_),
    .Y(_00112_));
 sky130_fd_sc_hd__clkinv_2 _19844_ (.A(_03107_),
    .Y(_00113_));
 sky130_fd_sc_hd__clkinv_2 _19845_ (.A(_03107_),
    .Y(_00114_));
 sky130_fd_sc_hd__clkinv_2 _19846_ (.A(_03107_),
    .Y(_00115_));
 sky130_fd_sc_hd__clkinv_2 _19847_ (.A(_03107_),
    .Y(_00116_));
 sky130_fd_sc_hd__buf_4 _19848_ (.A(_02862_),
    .X(_03108_));
 sky130_fd_sc_hd__clkinv_2 _19849_ (.A(_03108_),
    .Y(_00117_));
 sky130_fd_sc_hd__clkinv_2 _19850_ (.A(_03108_),
    .Y(_00118_));
 sky130_fd_sc_hd__clkinv_2 _19851_ (.A(_03108_),
    .Y(_00119_));
 sky130_fd_sc_hd__clkinv_2 _19852_ (.A(_03108_),
    .Y(_00120_));
 sky130_fd_sc_hd__clkinv_2 _19853_ (.A(_03108_),
    .Y(_00121_));
 sky130_fd_sc_hd__clkinv_2 _19854_ (.A(_03108_),
    .Y(_00122_));
 sky130_fd_sc_hd__clkinv_2 _19855_ (.A(_03108_),
    .Y(_00123_));
 sky130_fd_sc_hd__clkinv_2 _19856_ (.A(_03108_),
    .Y(_00124_));
 sky130_fd_sc_hd__clkinv_2 _19857_ (.A(_03108_),
    .Y(_00125_));
 sky130_fd_sc_hd__clkinv_2 _19858_ (.A(_03108_),
    .Y(_00126_));
 sky130_fd_sc_hd__buf_4 _19859_ (.A(_02862_),
    .X(_03109_));
 sky130_fd_sc_hd__clkinv_2 _19860_ (.A(_03109_),
    .Y(_00127_));
 sky130_fd_sc_hd__clkinv_2 _19861_ (.A(_03109_),
    .Y(_00128_));
 sky130_fd_sc_hd__clkinv_2 _19862_ (.A(_03109_),
    .Y(_00129_));
 sky130_fd_sc_hd__clkinv_2 _19863_ (.A(_03109_),
    .Y(_00130_));
 sky130_fd_sc_hd__clkinv_2 _19864_ (.A(_03109_),
    .Y(_00131_));
 sky130_fd_sc_hd__clkinv_2 _19865_ (.A(_03109_),
    .Y(_00132_));
 sky130_fd_sc_hd__clkinv_2 _19866_ (.A(_03109_),
    .Y(_00133_));
 sky130_fd_sc_hd__clkinv_2 _19867_ (.A(_03109_),
    .Y(_00134_));
 sky130_fd_sc_hd__clkinv_2 _19868_ (.A(_03109_),
    .Y(_00135_));
 sky130_fd_sc_hd__clkinv_2 _19869_ (.A(_03109_),
    .Y(_00136_));
 sky130_fd_sc_hd__buf_4 _19870_ (.A(_02862_),
    .X(_03110_));
 sky130_fd_sc_hd__clkinv_2 _19871_ (.A(_03110_),
    .Y(_00137_));
 sky130_fd_sc_hd__clkinv_2 _19872_ (.A(_03110_),
    .Y(_00138_));
 sky130_fd_sc_hd__clkinv_2 _19873_ (.A(_03110_),
    .Y(_00139_));
 sky130_fd_sc_hd__clkinv_2 _19874_ (.A(_03110_),
    .Y(_00140_));
 sky130_fd_sc_hd__clkinv_2 _19875_ (.A(_03110_),
    .Y(_00141_));
 sky130_fd_sc_hd__clkinv_2 _19876_ (.A(_03110_),
    .Y(_00142_));
 sky130_fd_sc_hd__clkinv_2 _19877_ (.A(_03110_),
    .Y(_00143_));
 sky130_fd_sc_hd__clkinv_2 _19878_ (.A(_03110_),
    .Y(_00144_));
 sky130_fd_sc_hd__clkinv_2 _19879_ (.A(_03110_),
    .Y(_00145_));
 sky130_fd_sc_hd__clkinv_2 _19880_ (.A(_03110_),
    .Y(_00146_));
 sky130_fd_sc_hd__buf_4 _19881_ (.A(_02862_),
    .X(_03111_));
 sky130_fd_sc_hd__clkinv_2 _19882_ (.A(_03111_),
    .Y(_00147_));
 sky130_fd_sc_hd__clkinv_2 _19883_ (.A(_03111_),
    .Y(_00148_));
 sky130_fd_sc_hd__clkinv_2 _19884_ (.A(_03111_),
    .Y(_00149_));
 sky130_fd_sc_hd__clkinv_2 _19885_ (.A(_03111_),
    .Y(_00150_));
 sky130_fd_sc_hd__clkinv_2 _19886_ (.A(_03111_),
    .Y(_00151_));
 sky130_fd_sc_hd__clkinv_2 _19887_ (.A(_03111_),
    .Y(_00152_));
 sky130_fd_sc_hd__clkinv_2 _19888_ (.A(_03111_),
    .Y(_00153_));
 sky130_fd_sc_hd__clkinv_2 _19889_ (.A(_03111_),
    .Y(_00154_));
 sky130_fd_sc_hd__clkinv_2 _19890_ (.A(_03111_),
    .Y(_00155_));
 sky130_fd_sc_hd__clkinv_2 _19891_ (.A(_03111_),
    .Y(_00156_));
 sky130_fd_sc_hd__buf_4 _19892_ (.A(_02862_),
    .X(_03112_));
 sky130_fd_sc_hd__clkinv_2 _19893_ (.A(_03112_),
    .Y(_00157_));
 sky130_fd_sc_hd__clkinv_2 _19894_ (.A(_03112_),
    .Y(_00158_));
 sky130_fd_sc_hd__clkinv_2 _19895_ (.A(_03112_),
    .Y(_00159_));
 sky130_fd_sc_hd__clkinv_2 _19896_ (.A(_03112_),
    .Y(_00160_));
 sky130_fd_sc_hd__clkinv_2 _19897_ (.A(_03112_),
    .Y(_00161_));
 sky130_fd_sc_hd__clkinv_2 _19898_ (.A(_03112_),
    .Y(_00162_));
 sky130_fd_sc_hd__clkinv_2 _19899_ (.A(_03112_),
    .Y(_00163_));
 sky130_fd_sc_hd__clkinv_2 _19900_ (.A(_03112_),
    .Y(_00164_));
 sky130_fd_sc_hd__clkinv_2 _19901_ (.A(_03112_),
    .Y(_00165_));
 sky130_fd_sc_hd__clkinv_2 _19902_ (.A(_03112_),
    .Y(_00166_));
 sky130_fd_sc_hd__buf_4 _19903_ (.A(_02862_),
    .X(_03113_));
 sky130_fd_sc_hd__clkinv_2 _19904_ (.A(_03113_),
    .Y(_00167_));
 sky130_fd_sc_hd__clkinv_2 _19905_ (.A(_03113_),
    .Y(_00168_));
 sky130_fd_sc_hd__clkinv_2 _19906_ (.A(_03113_),
    .Y(_00169_));
 sky130_fd_sc_hd__clkinv_2 _19907_ (.A(_03113_),
    .Y(_00170_));
 sky130_fd_sc_hd__clkinv_2 _19908_ (.A(_03113_),
    .Y(_00171_));
 sky130_fd_sc_hd__clkinv_2 _19909_ (.A(_03113_),
    .Y(_00172_));
 sky130_fd_sc_hd__clkinv_2 _19910_ (.A(_03113_),
    .Y(_00173_));
 sky130_fd_sc_hd__clkinv_2 _19911_ (.A(_03113_),
    .Y(_00174_));
 sky130_fd_sc_hd__clkinv_2 _19912_ (.A(_03113_),
    .Y(_00175_));
 sky130_fd_sc_hd__clkinv_2 _19913_ (.A(_03113_),
    .Y(_00176_));
 sky130_fd_sc_hd__buf_4 _19914_ (.A(_04702_),
    .X(_03114_));
 sky130_fd_sc_hd__buf_4 _19915_ (.A(_03114_),
    .X(_03115_));
 sky130_fd_sc_hd__clkinv_2 _19916_ (.A(_03115_),
    .Y(_00177_));
 sky130_fd_sc_hd__clkinv_2 _19917_ (.A(_03115_),
    .Y(_00178_));
 sky130_fd_sc_hd__clkinv_2 _19918_ (.A(_03115_),
    .Y(_00179_));
 sky130_fd_sc_hd__clkinv_2 _19919_ (.A(_03115_),
    .Y(_00180_));
 sky130_fd_sc_hd__clkinv_2 _19920_ (.A(_03115_),
    .Y(_00181_));
 sky130_fd_sc_hd__clkinv_2 _19921_ (.A(_03115_),
    .Y(_00182_));
 sky130_fd_sc_hd__clkinv_2 _19922_ (.A(_03115_),
    .Y(_00183_));
 sky130_fd_sc_hd__clkinv_2 _19923_ (.A(_03115_),
    .Y(_00184_));
 sky130_fd_sc_hd__clkinv_2 _19924_ (.A(_03115_),
    .Y(_00185_));
 sky130_fd_sc_hd__clkinv_2 _19925_ (.A(_03115_),
    .Y(_00186_));
 sky130_fd_sc_hd__buf_4 _19926_ (.A(_03114_),
    .X(_03116_));
 sky130_fd_sc_hd__clkinv_2 _19927_ (.A(_03116_),
    .Y(_00187_));
 sky130_fd_sc_hd__clkinv_2 _19928_ (.A(_03116_),
    .Y(_00188_));
 sky130_fd_sc_hd__clkinv_2 _19929_ (.A(_03116_),
    .Y(_00189_));
 sky130_fd_sc_hd__clkinv_2 _19930_ (.A(_03116_),
    .Y(_00190_));
 sky130_fd_sc_hd__clkinv_2 _19931_ (.A(_03116_),
    .Y(_00191_));
 sky130_fd_sc_hd__clkinv_2 _19932_ (.A(_03116_),
    .Y(_00192_));
 sky130_fd_sc_hd__clkinv_2 _19933_ (.A(_03116_),
    .Y(_00193_));
 sky130_fd_sc_hd__clkinv_2 _19934_ (.A(_03116_),
    .Y(_00194_));
 sky130_fd_sc_hd__clkinv_2 _19935_ (.A(_03116_),
    .Y(_00195_));
 sky130_fd_sc_hd__clkinv_2 _19936_ (.A(_03116_),
    .Y(_00196_));
 sky130_fd_sc_hd__buf_4 _19937_ (.A(_03114_),
    .X(_03117_));
 sky130_fd_sc_hd__clkinv_2 _19938_ (.A(_03117_),
    .Y(_00197_));
 sky130_fd_sc_hd__clkinv_2 _19939_ (.A(_03117_),
    .Y(_00198_));
 sky130_fd_sc_hd__clkinv_2 _19940_ (.A(_03117_),
    .Y(_00199_));
 sky130_fd_sc_hd__clkinv_2 _19941_ (.A(_03117_),
    .Y(_00200_));
 sky130_fd_sc_hd__clkinv_2 _19942_ (.A(_03117_),
    .Y(_00201_));
 sky130_fd_sc_hd__clkinv_2 _19943_ (.A(_03117_),
    .Y(_00202_));
 sky130_fd_sc_hd__clkinv_2 _19944_ (.A(_03117_),
    .Y(_00203_));
 sky130_fd_sc_hd__clkinv_2 _19945_ (.A(_03117_),
    .Y(_00204_));
 sky130_fd_sc_hd__clkinv_2 _19946_ (.A(_03117_),
    .Y(_00205_));
 sky130_fd_sc_hd__clkinv_2 _19947_ (.A(_03117_),
    .Y(_00206_));
 sky130_fd_sc_hd__buf_4 _19948_ (.A(_03114_),
    .X(_03118_));
 sky130_fd_sc_hd__clkinv_2 _19949_ (.A(_03118_),
    .Y(_00207_));
 sky130_fd_sc_hd__clkinv_2 _19950_ (.A(_03118_),
    .Y(_00208_));
 sky130_fd_sc_hd__clkinv_2 _19951_ (.A(_03118_),
    .Y(_00209_));
 sky130_fd_sc_hd__clkinv_2 _19952_ (.A(_03118_),
    .Y(_00210_));
 sky130_fd_sc_hd__clkinv_2 _19953_ (.A(_03118_),
    .Y(_00211_));
 sky130_fd_sc_hd__clkinv_2 _19954_ (.A(_03118_),
    .Y(_00212_));
 sky130_fd_sc_hd__clkinv_2 _19955_ (.A(_03118_),
    .Y(_00213_));
 sky130_fd_sc_hd__clkinv_2 _19956_ (.A(_03118_),
    .Y(_00214_));
 sky130_fd_sc_hd__clkinv_2 _19957_ (.A(_03118_),
    .Y(_00215_));
 sky130_fd_sc_hd__clkinv_2 _19958_ (.A(_03118_),
    .Y(_00216_));
 sky130_fd_sc_hd__clkbuf_8 _19959_ (.A(_03114_),
    .X(_03119_));
 sky130_fd_sc_hd__clkinv_2 _19960_ (.A(_03119_),
    .Y(_00217_));
 sky130_fd_sc_hd__clkinv_2 _19961_ (.A(_03119_),
    .Y(_00218_));
 sky130_fd_sc_hd__clkinv_2 _19962_ (.A(_03119_),
    .Y(_00219_));
 sky130_fd_sc_hd__clkinv_2 _19963_ (.A(_03119_),
    .Y(_00220_));
 sky130_fd_sc_hd__clkinv_2 _19964_ (.A(_03119_),
    .Y(_00221_));
 sky130_fd_sc_hd__clkinv_2 _19965_ (.A(_03119_),
    .Y(_00222_));
 sky130_fd_sc_hd__clkinv_2 _19966_ (.A(_03119_),
    .Y(_00223_));
 sky130_fd_sc_hd__clkinv_2 _19967_ (.A(_03119_),
    .Y(_00224_));
 sky130_fd_sc_hd__clkinv_2 _19968_ (.A(_03119_),
    .Y(_00225_));
 sky130_fd_sc_hd__clkinv_2 _19969_ (.A(_03119_),
    .Y(_00226_));
 sky130_fd_sc_hd__clkbuf_8 _19970_ (.A(_03114_),
    .X(_03120_));
 sky130_fd_sc_hd__clkinv_2 _19971_ (.A(_03120_),
    .Y(_00227_));
 sky130_fd_sc_hd__clkinv_2 _19972_ (.A(_03120_),
    .Y(_00228_));
 sky130_fd_sc_hd__clkinv_2 _19973_ (.A(_03120_),
    .Y(_00229_));
 sky130_fd_sc_hd__clkinv_2 _19974_ (.A(_03120_),
    .Y(_00230_));
 sky130_fd_sc_hd__clkinv_2 _19975_ (.A(_03120_),
    .Y(_00231_));
 sky130_fd_sc_hd__clkinv_2 _19976_ (.A(_03120_),
    .Y(_00232_));
 sky130_fd_sc_hd__clkinv_2 _19977_ (.A(_03120_),
    .Y(_00233_));
 sky130_fd_sc_hd__clkinv_2 _19978_ (.A(_03120_),
    .Y(_00234_));
 sky130_fd_sc_hd__clkinv_2 _19979_ (.A(_03120_),
    .Y(_00235_));
 sky130_fd_sc_hd__clkinv_2 _19980_ (.A(_03120_),
    .Y(_00236_));
 sky130_fd_sc_hd__buf_4 _19981_ (.A(_03114_),
    .X(_03121_));
 sky130_fd_sc_hd__clkinv_2 _19982_ (.A(_03121_),
    .Y(_00237_));
 sky130_fd_sc_hd__clkinv_2 _19983_ (.A(_03121_),
    .Y(_00238_));
 sky130_fd_sc_hd__clkinv_2 _19984_ (.A(_03121_),
    .Y(_00239_));
 sky130_fd_sc_hd__clkinv_2 _19985_ (.A(_03121_),
    .Y(_00240_));
 sky130_fd_sc_hd__clkinv_2 _19986_ (.A(_03121_),
    .Y(_00241_));
 sky130_fd_sc_hd__clkinv_2 _19987_ (.A(_03121_),
    .Y(_00242_));
 sky130_fd_sc_hd__clkinv_2 _19988_ (.A(_03121_),
    .Y(_00243_));
 sky130_fd_sc_hd__clkinv_2 _19989_ (.A(_03121_),
    .Y(_00244_));
 sky130_fd_sc_hd__clkinv_2 _19990_ (.A(_03121_),
    .Y(_00245_));
 sky130_fd_sc_hd__clkinv_2 _19991_ (.A(_03121_),
    .Y(_00246_));
 sky130_fd_sc_hd__buf_4 _19992_ (.A(_03114_),
    .X(_03122_));
 sky130_fd_sc_hd__clkinv_2 _19993_ (.A(_03122_),
    .Y(_00247_));
 sky130_fd_sc_hd__clkinv_2 _19994_ (.A(_03122_),
    .Y(_00248_));
 sky130_fd_sc_hd__clkinv_2 _19995_ (.A(_03122_),
    .Y(_00249_));
 sky130_fd_sc_hd__clkinv_2 _19996_ (.A(_03122_),
    .Y(_00250_));
 sky130_fd_sc_hd__clkinv_2 _19997_ (.A(_03122_),
    .Y(_00251_));
 sky130_fd_sc_hd__clkinv_2 _19998_ (.A(_03122_),
    .Y(_00252_));
 sky130_fd_sc_hd__clkinv_2 _19999_ (.A(_03122_),
    .Y(_00253_));
 sky130_fd_sc_hd__clkinv_2 _20000_ (.A(_03122_),
    .Y(_00254_));
 sky130_fd_sc_hd__clkinv_2 _20001_ (.A(_03122_),
    .Y(_00255_));
 sky130_fd_sc_hd__clkinv_2 _20002_ (.A(_03122_),
    .Y(_00256_));
 sky130_fd_sc_hd__buf_4 _20003_ (.A(_03114_),
    .X(_03123_));
 sky130_fd_sc_hd__clkinv_2 _20004_ (.A(_03123_),
    .Y(_00257_));
 sky130_fd_sc_hd__clkinv_2 _20005_ (.A(_03123_),
    .Y(_00258_));
 sky130_fd_sc_hd__clkinv_2 _20006_ (.A(_03123_),
    .Y(_00259_));
 sky130_fd_sc_hd__clkinv_2 _20007_ (.A(_03123_),
    .Y(_00260_));
 sky130_fd_sc_hd__clkinv_2 _20008_ (.A(_03123_),
    .Y(_00261_));
 sky130_fd_sc_hd__clkinv_2 _20009_ (.A(_03123_),
    .Y(_00262_));
 sky130_fd_sc_hd__clkinv_2 _20010_ (.A(_03123_),
    .Y(_00263_));
 sky130_fd_sc_hd__clkinv_2 _20011_ (.A(_03123_),
    .Y(_00264_));
 sky130_fd_sc_hd__clkinv_2 _20012_ (.A(_03123_),
    .Y(_00265_));
 sky130_fd_sc_hd__clkinv_2 _20013_ (.A(_03123_),
    .Y(_00266_));
 sky130_fd_sc_hd__buf_4 _20014_ (.A(_03114_),
    .X(_03124_));
 sky130_fd_sc_hd__clkinv_2 _20015_ (.A(_03124_),
    .Y(_00267_));
 sky130_fd_sc_hd__clkinv_2 _20016_ (.A(_03124_),
    .Y(_00268_));
 sky130_fd_sc_hd__clkinv_2 _20017_ (.A(_03124_),
    .Y(_00269_));
 sky130_fd_sc_hd__clkinv_2 _20018_ (.A(_03124_),
    .Y(_00270_));
 sky130_fd_sc_hd__clkinv_2 _20019_ (.A(_03124_),
    .Y(_00271_));
 sky130_fd_sc_hd__clkinv_2 _20020_ (.A(_03124_),
    .Y(_00272_));
 sky130_fd_sc_hd__clkinv_2 _20021_ (.A(_03124_),
    .Y(_00273_));
 sky130_fd_sc_hd__clkinv_2 _20022_ (.A(_03124_),
    .Y(_00274_));
 sky130_fd_sc_hd__clkinv_2 _20023_ (.A(_03124_),
    .Y(_00275_));
 sky130_fd_sc_hd__clkinv_2 _20024_ (.A(_03124_),
    .Y(_00276_));
 sky130_fd_sc_hd__buf_4 _20025_ (.A(_04702_),
    .X(_03125_));
 sky130_fd_sc_hd__buf_4 _20026_ (.A(_03125_),
    .X(_03126_));
 sky130_fd_sc_hd__clkinv_2 _20027_ (.A(_03126_),
    .Y(_00277_));
 sky130_fd_sc_hd__clkinv_2 _20028_ (.A(_03126_),
    .Y(_00278_));
 sky130_fd_sc_hd__clkinv_2 _20029_ (.A(_03126_),
    .Y(_00279_));
 sky130_fd_sc_hd__clkinv_2 _20030_ (.A(_03126_),
    .Y(_00280_));
 sky130_fd_sc_hd__clkinv_2 _20031_ (.A(_03126_),
    .Y(_00281_));
 sky130_fd_sc_hd__clkinv_2 _20032_ (.A(_03126_),
    .Y(_00282_));
 sky130_fd_sc_hd__clkinv_2 _20033_ (.A(_03126_),
    .Y(_00283_));
 sky130_fd_sc_hd__clkinv_2 _20034_ (.A(_03126_),
    .Y(_00284_));
 sky130_fd_sc_hd__clkinv_2 _20035_ (.A(_03126_),
    .Y(_00285_));
 sky130_fd_sc_hd__clkinv_2 _20036_ (.A(_03126_),
    .Y(_00286_));
 sky130_fd_sc_hd__clkbuf_8 _20037_ (.A(_03125_),
    .X(_03127_));
 sky130_fd_sc_hd__clkinv_2 _20038_ (.A(_03127_),
    .Y(_00287_));
 sky130_fd_sc_hd__clkinv_2 _20039_ (.A(_03127_),
    .Y(_00288_));
 sky130_fd_sc_hd__clkinv_2 _20040_ (.A(_03127_),
    .Y(_00289_));
 sky130_fd_sc_hd__clkinv_2 _20041_ (.A(_03127_),
    .Y(_00290_));
 sky130_fd_sc_hd__clkinv_2 _20042_ (.A(_03127_),
    .Y(_00291_));
 sky130_fd_sc_hd__clkinv_2 _20043_ (.A(_03127_),
    .Y(_00292_));
 sky130_fd_sc_hd__clkinv_2 _20044_ (.A(_03127_),
    .Y(_00293_));
 sky130_fd_sc_hd__clkinv_2 _20045_ (.A(_03127_),
    .Y(_00294_));
 sky130_fd_sc_hd__clkinv_2 _20046_ (.A(_03127_),
    .Y(_00295_));
 sky130_fd_sc_hd__clkinv_2 _20047_ (.A(_03127_),
    .Y(_00296_));
 sky130_fd_sc_hd__buf_4 _20048_ (.A(_03125_),
    .X(_03128_));
 sky130_fd_sc_hd__clkinv_2 _20049_ (.A(_03128_),
    .Y(_00297_));
 sky130_fd_sc_hd__clkinv_2 _20050_ (.A(_03128_),
    .Y(_00298_));
 sky130_fd_sc_hd__clkinv_2 _20051_ (.A(_03128_),
    .Y(_00299_));
 sky130_fd_sc_hd__clkinv_2 _20052_ (.A(_03128_),
    .Y(_00300_));
 sky130_fd_sc_hd__clkinv_2 _20053_ (.A(_03128_),
    .Y(_00301_));
 sky130_fd_sc_hd__clkinv_2 _20054_ (.A(_03128_),
    .Y(_00302_));
 sky130_fd_sc_hd__clkinv_2 _20055_ (.A(_03128_),
    .Y(_00303_));
 sky130_fd_sc_hd__clkinv_2 _20056_ (.A(_03128_),
    .Y(_00304_));
 sky130_fd_sc_hd__clkinv_2 _20057_ (.A(_03128_),
    .Y(_00305_));
 sky130_fd_sc_hd__clkinv_2 _20058_ (.A(_03128_),
    .Y(_00306_));
 sky130_fd_sc_hd__buf_4 _20059_ (.A(_03125_),
    .X(_03129_));
 sky130_fd_sc_hd__clkinv_2 _20060_ (.A(_03129_),
    .Y(_00307_));
 sky130_fd_sc_hd__clkinv_2 _20061_ (.A(_03129_),
    .Y(_00308_));
 sky130_fd_sc_hd__clkinv_2 _20062_ (.A(_03129_),
    .Y(_00309_));
 sky130_fd_sc_hd__clkinv_2 _20063_ (.A(_03129_),
    .Y(_00310_));
 sky130_fd_sc_hd__clkinv_2 _20064_ (.A(_03129_),
    .Y(_00311_));
 sky130_fd_sc_hd__clkinv_2 _20065_ (.A(_03129_),
    .Y(_00312_));
 sky130_fd_sc_hd__clkinv_2 _20066_ (.A(_03129_),
    .Y(_00313_));
 sky130_fd_sc_hd__clkinv_2 _20067_ (.A(_03129_),
    .Y(_00314_));
 sky130_fd_sc_hd__clkinv_2 _20068_ (.A(_03129_),
    .Y(_00315_));
 sky130_fd_sc_hd__clkinv_2 _20069_ (.A(_03129_),
    .Y(_00316_));
 sky130_fd_sc_hd__buf_6 _20070_ (.A(_03125_),
    .X(_03130_));
 sky130_fd_sc_hd__clkinv_2 _20071_ (.A(_03130_),
    .Y(_00317_));
 sky130_fd_sc_hd__clkinv_2 _20072_ (.A(_03130_),
    .Y(_00318_));
 sky130_fd_sc_hd__clkinv_2 _20073_ (.A(_03130_),
    .Y(_00319_));
 sky130_fd_sc_hd__clkinv_2 _20074_ (.A(_03130_),
    .Y(_00320_));
 sky130_fd_sc_hd__clkinv_2 _20075_ (.A(_03130_),
    .Y(_00321_));
 sky130_fd_sc_hd__clkinv_2 _20076_ (.A(_03130_),
    .Y(_00322_));
 sky130_fd_sc_hd__clkinv_2 _20077_ (.A(_03130_),
    .Y(_00323_));
 sky130_fd_sc_hd__clkinv_2 _20078_ (.A(_03130_),
    .Y(_00324_));
 sky130_fd_sc_hd__clkinv_2 _20079_ (.A(_03130_),
    .Y(_00325_));
 sky130_fd_sc_hd__clkinv_2 _20080_ (.A(_03130_),
    .Y(_00326_));
 sky130_fd_sc_hd__buf_4 _20081_ (.A(_03125_),
    .X(_03131_));
 sky130_fd_sc_hd__clkinv_2 _20082_ (.A(_03131_),
    .Y(_00327_));
 sky130_fd_sc_hd__clkinv_2 _20083_ (.A(_03131_),
    .Y(_00328_));
 sky130_fd_sc_hd__clkinv_2 _20084_ (.A(_03131_),
    .Y(_00329_));
 sky130_fd_sc_hd__clkinv_2 _20085_ (.A(_03131_),
    .Y(_00330_));
 sky130_fd_sc_hd__clkinv_2 _20086_ (.A(_03131_),
    .Y(_00331_));
 sky130_fd_sc_hd__clkinv_2 _20087_ (.A(_03131_),
    .Y(_00332_));
 sky130_fd_sc_hd__clkinv_2 _20088_ (.A(_03131_),
    .Y(_00333_));
 sky130_fd_sc_hd__clkinv_2 _20089_ (.A(_03131_),
    .Y(_00334_));
 sky130_fd_sc_hd__clkinv_2 _20090_ (.A(_03131_),
    .Y(_00335_));
 sky130_fd_sc_hd__clkinv_2 _20091_ (.A(_03131_),
    .Y(_00336_));
 sky130_fd_sc_hd__nor2_1 _20092_ (.A(\gpout5.clk_div[0] ),
    .B(_03003_),
    .Y(_01304_));
 sky130_fd_sc_hd__nand2_1 _20093_ (.A(\gpout5.clk_div[1] ),
    .B(\gpout5.clk_div[0] ),
    .Y(_03132_));
 sky130_fd_sc_hd__or2_1 _20094_ (.A(\gpout5.clk_div[1] ),
    .B(\gpout5.clk_div[0] ),
    .X(_03133_));
 sky130_fd_sc_hd__and3_1 _20095_ (.A(_09247_),
    .B(_03132_),
    .C(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__clkbuf_1 _20096_ (.A(_03134_),
    .X(_01305_));
 sky130_fd_sc_hd__nand2_1 _20097_ (.A(\rbzero.traced_texa[-12] ),
    .B(\rbzero.texV[-12] ),
    .Y(_03135_));
 sky130_fd_sc_hd__or2_1 _20098_ (.A(\rbzero.traced_texa[-12] ),
    .B(\rbzero.texV[-12] ),
    .X(_03136_));
 sky130_fd_sc_hd__clkbuf_4 _20099_ (.A(_02708_),
    .X(_03137_));
 sky130_fd_sc_hd__a32o_1 _20100_ (.A1(_03093_),
    .A2(_03135_),
    .A3(_03136_),
    .B1(_03137_),
    .B2(\rbzero.texV[-12] ),
    .X(_01306_));
 sky130_fd_sc_hd__or2_1 _20101_ (.A(\rbzero.traced_texa[-11] ),
    .B(\rbzero.texV[-11] ),
    .X(_03138_));
 sky130_fd_sc_hd__nand2_1 _20102_ (.A(\rbzero.traced_texa[-11] ),
    .B(\rbzero.texV[-11] ),
    .Y(_03139_));
 sky130_fd_sc_hd__nand3b_1 _20103_ (.A_N(_03135_),
    .B(_03138_),
    .C(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hd__a21bo_1 _20104_ (.A1(_03138_),
    .A2(_03139_),
    .B1_N(_03135_),
    .X(_03141_));
 sky130_fd_sc_hd__a32o_1 _20105_ (.A1(_03093_),
    .A2(_03140_),
    .A3(_03141_),
    .B1(_03137_),
    .B2(\rbzero.texV[-11] ),
    .X(_01307_));
 sky130_fd_sc_hd__buf_2 _20106_ (.A(_09245_),
    .X(_03142_));
 sky130_fd_sc_hd__and2_1 _20107_ (.A(_03139_),
    .B(_03140_),
    .X(_03143_));
 sky130_fd_sc_hd__nor2_1 _20108_ (.A(\rbzero.traced_texa[-10] ),
    .B(\rbzero.texV[-10] ),
    .Y(_03144_));
 sky130_fd_sc_hd__nand2_1 _20109_ (.A(\rbzero.traced_texa[-10] ),
    .B(\rbzero.texV[-10] ),
    .Y(_03145_));
 sky130_fd_sc_hd__and2b_1 _20110_ (.A_N(_03144_),
    .B(_03145_),
    .X(_03146_));
 sky130_fd_sc_hd__xnor2_1 _20111_ (.A(_03143_),
    .B(_03146_),
    .Y(_03147_));
 sky130_fd_sc_hd__a22o_1 _20112_ (.A1(\rbzero.texV[-10] ),
    .A2(_02989_),
    .B1(_03142_),
    .B2(_03147_),
    .X(_01308_));
 sky130_fd_sc_hd__or2_1 _20113_ (.A(\rbzero.traced_texa[-9] ),
    .B(\rbzero.texV[-9] ),
    .X(_03148_));
 sky130_fd_sc_hd__nand2_1 _20114_ (.A(\rbzero.traced_texa[-9] ),
    .B(\rbzero.texV[-9] ),
    .Y(_03149_));
 sky130_fd_sc_hd__nand2_1 _20115_ (.A(_03148_),
    .B(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hd__o21ai_1 _20116_ (.A1(_03143_),
    .A2(_03144_),
    .B1(_03145_),
    .Y(_03151_));
 sky130_fd_sc_hd__xnor2_1 _20117_ (.A(_03150_),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__a22o_1 _20118_ (.A1(\rbzero.texV[-9] ),
    .A2(_02989_),
    .B1(_03142_),
    .B2(_03152_),
    .X(_01309_));
 sky130_fd_sc_hd__nor2_1 _20119_ (.A(\rbzero.traced_texa[-8] ),
    .B(\rbzero.texV[-8] ),
    .Y(_03153_));
 sky130_fd_sc_hd__and2_1 _20120_ (.A(\rbzero.traced_texa[-8] ),
    .B(\rbzero.texV[-8] ),
    .X(_03154_));
 sky130_fd_sc_hd__a21boi_1 _20121_ (.A1(_03148_),
    .A2(_03151_),
    .B1_N(_03149_),
    .Y(_03155_));
 sky130_fd_sc_hd__o21ai_1 _20122_ (.A1(_03153_),
    .A2(_03154_),
    .B1(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__or3_1 _20123_ (.A(_03153_),
    .B(_03154_),
    .C(_03155_),
    .X(_03157_));
 sky130_fd_sc_hd__a32o_1 _20124_ (.A1(_03093_),
    .A2(_03156_),
    .A3(_03157_),
    .B1(_03137_),
    .B2(\rbzero.texV[-8] ),
    .X(_01310_));
 sky130_fd_sc_hd__or2_1 _20125_ (.A(\rbzero.traced_texa[-7] ),
    .B(\rbzero.texV[-7] ),
    .X(_03158_));
 sky130_fd_sc_hd__nand2_1 _20126_ (.A(\rbzero.traced_texa[-7] ),
    .B(\rbzero.texV[-7] ),
    .Y(_03159_));
 sky130_fd_sc_hd__o21bai_1 _20127_ (.A1(_03153_),
    .A2(_03155_),
    .B1_N(_03154_),
    .Y(_03160_));
 sky130_fd_sc_hd__nand3_1 _20128_ (.A(_03158_),
    .B(_03159_),
    .C(_03160_),
    .Y(_03161_));
 sky130_fd_sc_hd__a21o_1 _20129_ (.A1(_03158_),
    .A2(_03159_),
    .B1(_03160_),
    .X(_03162_));
 sky130_fd_sc_hd__a32o_1 _20130_ (.A1(_03093_),
    .A2(_03161_),
    .A3(_03162_),
    .B1(_03137_),
    .B2(\rbzero.texV[-7] ),
    .X(_01311_));
 sky130_fd_sc_hd__nor2_1 _20131_ (.A(\rbzero.traced_texa[-6] ),
    .B(\rbzero.texV[-6] ),
    .Y(_03163_));
 sky130_fd_sc_hd__and2_1 _20132_ (.A(\rbzero.traced_texa[-6] ),
    .B(\rbzero.texV[-6] ),
    .X(_03164_));
 sky130_fd_sc_hd__a21boi_1 _20133_ (.A1(_03158_),
    .A2(_03160_),
    .B1_N(_03159_),
    .Y(_03165_));
 sky130_fd_sc_hd__or3_1 _20134_ (.A(_03163_),
    .B(_03164_),
    .C(_03165_),
    .X(_03166_));
 sky130_fd_sc_hd__o21ai_1 _20135_ (.A1(_03163_),
    .A2(_03164_),
    .B1(_03165_),
    .Y(_03167_));
 sky130_fd_sc_hd__a32o_1 _20136_ (.A1(_03093_),
    .A2(_03166_),
    .A3(_03167_),
    .B1(_03137_),
    .B2(\rbzero.texV[-6] ),
    .X(_01312_));
 sky130_fd_sc_hd__xnor2_1 _20137_ (.A(\rbzero.traced_texa[-5] ),
    .B(\rbzero.texV[-5] ),
    .Y(_03168_));
 sky130_fd_sc_hd__o21bai_1 _20138_ (.A1(_03163_),
    .A2(_03165_),
    .B1_N(_03164_),
    .Y(_03169_));
 sky130_fd_sc_hd__xnor2_1 _20139_ (.A(_03168_),
    .B(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__a22o_1 _20140_ (.A1(\rbzero.texV[-5] ),
    .A2(_02989_),
    .B1(_03142_),
    .B2(_03170_),
    .X(_01313_));
 sky130_fd_sc_hd__nor2_1 _20141_ (.A(\rbzero.traced_texa[-4] ),
    .B(\rbzero.texV[-4] ),
    .Y(_03171_));
 sky130_fd_sc_hd__nand2_1 _20142_ (.A(\rbzero.traced_texa[-4] ),
    .B(\rbzero.texV[-4] ),
    .Y(_03172_));
 sky130_fd_sc_hd__and2b_1 _20143_ (.A_N(_03171_),
    .B(_03172_),
    .X(_03173_));
 sky130_fd_sc_hd__a21o_1 _20144_ (.A1(\rbzero.traced_texa[-5] ),
    .A2(\rbzero.texV[-5] ),
    .B1(_03169_),
    .X(_03174_));
 sky130_fd_sc_hd__o21ai_1 _20145_ (.A1(\rbzero.traced_texa[-5] ),
    .A2(\rbzero.texV[-5] ),
    .B1(_03174_),
    .Y(_03175_));
 sky130_fd_sc_hd__xnor2_1 _20146_ (.A(_03173_),
    .B(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__a22o_1 _20147_ (.A1(\rbzero.texV[-4] ),
    .A2(_02989_),
    .B1(_03142_),
    .B2(_03176_),
    .X(_01314_));
 sky130_fd_sc_hd__or2_1 _20148_ (.A(\rbzero.traced_texa[-3] ),
    .B(\rbzero.texV[-3] ),
    .X(_03177_));
 sky130_fd_sc_hd__nand2_1 _20149_ (.A(\rbzero.traced_texa[-3] ),
    .B(\rbzero.texV[-3] ),
    .Y(_03178_));
 sky130_fd_sc_hd__o21ai_1 _20150_ (.A1(_03171_),
    .A2(_03175_),
    .B1(_03172_),
    .Y(_03179_));
 sky130_fd_sc_hd__a21o_1 _20151_ (.A1(_03177_),
    .A2(_03178_),
    .B1(_03179_),
    .X(_03180_));
 sky130_fd_sc_hd__nand3_1 _20152_ (.A(_03177_),
    .B(_03178_),
    .C(_03179_),
    .Y(_03181_));
 sky130_fd_sc_hd__a32o_1 _20153_ (.A1(_03093_),
    .A2(_03180_),
    .A3(_03181_),
    .B1(_03064_),
    .B2(\rbzero.texV[-3] ),
    .X(_01315_));
 sky130_fd_sc_hd__nor2_1 _20154_ (.A(\rbzero.traced_texa[-2] ),
    .B(\rbzero.texV[-2] ),
    .Y(_03182_));
 sky130_fd_sc_hd__and2_1 _20155_ (.A(\rbzero.traced_texa[-2] ),
    .B(\rbzero.texV[-2] ),
    .X(_03183_));
 sky130_fd_sc_hd__or2_1 _20156_ (.A(_03182_),
    .B(_03183_),
    .X(_03184_));
 sky130_fd_sc_hd__a21boi_1 _20157_ (.A1(_03177_),
    .A2(_03179_),
    .B1_N(_03178_),
    .Y(_03185_));
 sky130_fd_sc_hd__xor2_1 _20158_ (.A(_03184_),
    .B(_03185_),
    .X(_03186_));
 sky130_fd_sc_hd__a22o_1 _20159_ (.A1(\rbzero.texV[-2] ),
    .A2(_02989_),
    .B1(_03142_),
    .B2(_03186_),
    .X(_01316_));
 sky130_fd_sc_hd__nor2_1 _20160_ (.A(_03184_),
    .B(_03185_),
    .Y(_03187_));
 sky130_fd_sc_hd__or2_1 _20161_ (.A(\rbzero.traced_texa[-1] ),
    .B(\rbzero.texV[-1] ),
    .X(_03188_));
 sky130_fd_sc_hd__nand2_1 _20162_ (.A(\rbzero.traced_texa[-1] ),
    .B(\rbzero.texV[-1] ),
    .Y(_03189_));
 sky130_fd_sc_hd__o211a_1 _20163_ (.A1(_03183_),
    .A2(_03187_),
    .B1(_03188_),
    .C1(_03189_),
    .X(_03190_));
 sky130_fd_sc_hd__inv_2 _20164_ (.A(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__a211o_1 _20165_ (.A1(_03188_),
    .A2(_03189_),
    .B1(_03183_),
    .C1(_03187_),
    .X(_03192_));
 sky130_fd_sc_hd__a32o_1 _20166_ (.A1(_03093_),
    .A2(_03191_),
    .A3(_03192_),
    .B1(_03064_),
    .B2(\rbzero.texV[-1] ),
    .X(_01317_));
 sky130_fd_sc_hd__or2_1 _20167_ (.A(\rbzero.traced_texa[0] ),
    .B(\rbzero.texV[0] ),
    .X(_03193_));
 sky130_fd_sc_hd__nand2_1 _20168_ (.A(\rbzero.traced_texa[0] ),
    .B(\rbzero.texV[0] ),
    .Y(_03194_));
 sky130_fd_sc_hd__nand2_1 _20169_ (.A(_03189_),
    .B(_03191_),
    .Y(_03195_));
 sky130_fd_sc_hd__a21o_1 _20170_ (.A1(_03193_),
    .A2(_03194_),
    .B1(_03195_),
    .X(_03196_));
 sky130_fd_sc_hd__and3_1 _20171_ (.A(_03193_),
    .B(_03194_),
    .C(_03195_),
    .X(_03197_));
 sky130_fd_sc_hd__inv_2 _20172_ (.A(_03197_),
    .Y(_03198_));
 sky130_fd_sc_hd__a32o_1 _20173_ (.A1(_03093_),
    .A2(_03196_),
    .A3(_03198_),
    .B1(_03064_),
    .B2(\rbzero.texV[0] ),
    .X(_01318_));
 sky130_fd_sc_hd__or2_1 _20174_ (.A(\rbzero.traced_texa[1] ),
    .B(\rbzero.texV[1] ),
    .X(_03199_));
 sky130_fd_sc_hd__nand2_1 _20175_ (.A(\rbzero.traced_texa[1] ),
    .B(\rbzero.texV[1] ),
    .Y(_03200_));
 sky130_fd_sc_hd__nand2_1 _20176_ (.A(_03194_),
    .B(_03198_),
    .Y(_03201_));
 sky130_fd_sc_hd__and3_1 _20177_ (.A(_03199_),
    .B(_03200_),
    .C(_03201_),
    .X(_03202_));
 sky130_fd_sc_hd__inv_2 _20178_ (.A(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__a21o_1 _20179_ (.A1(_03199_),
    .A2(_03200_),
    .B1(_03201_),
    .X(_03204_));
 sky130_fd_sc_hd__a32o_1 _20180_ (.A1(_03093_),
    .A2(_03203_),
    .A3(_03204_),
    .B1(_03064_),
    .B2(\rbzero.texV[1] ),
    .X(_01319_));
 sky130_fd_sc_hd__or2_1 _20181_ (.A(\rbzero.traced_texa[2] ),
    .B(\rbzero.texV[2] ),
    .X(_03205_));
 sky130_fd_sc_hd__nand2_1 _20182_ (.A(\rbzero.traced_texa[2] ),
    .B(\rbzero.texV[2] ),
    .Y(_03206_));
 sky130_fd_sc_hd__nand2_1 _20183_ (.A(_03200_),
    .B(_03203_),
    .Y(_03207_));
 sky130_fd_sc_hd__a21o_1 _20184_ (.A1(_03205_),
    .A2(_03206_),
    .B1(_03207_),
    .X(_03208_));
 sky130_fd_sc_hd__and3_1 _20185_ (.A(_03205_),
    .B(_03206_),
    .C(_03207_),
    .X(_03209_));
 sky130_fd_sc_hd__inv_2 _20186_ (.A(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__a32o_1 _20187_ (.A1(_09245_),
    .A2(_03208_),
    .A3(_03210_),
    .B1(_03064_),
    .B2(\rbzero.texV[2] ),
    .X(_01320_));
 sky130_fd_sc_hd__or2_1 _20188_ (.A(\rbzero.traced_texa[3] ),
    .B(\rbzero.texV[3] ),
    .X(_03211_));
 sky130_fd_sc_hd__nand2_1 _20189_ (.A(\rbzero.traced_texa[3] ),
    .B(\rbzero.texV[3] ),
    .Y(_03212_));
 sky130_fd_sc_hd__nand2_1 _20190_ (.A(_03206_),
    .B(_03210_),
    .Y(_03213_));
 sky130_fd_sc_hd__nand3_1 _20191_ (.A(_03211_),
    .B(_03212_),
    .C(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__a21o_1 _20192_ (.A1(_03211_),
    .A2(_03212_),
    .B1(_03213_),
    .X(_03215_));
 sky130_fd_sc_hd__a32o_1 _20193_ (.A1(_09245_),
    .A2(_03214_),
    .A3(_03215_),
    .B1(_03064_),
    .B2(\rbzero.texV[3] ),
    .X(_01321_));
 sky130_fd_sc_hd__a21boi_1 _20194_ (.A1(_03211_),
    .A2(_03213_),
    .B1_N(_03212_),
    .Y(_03216_));
 sky130_fd_sc_hd__nor2_1 _20195_ (.A(\rbzero.traced_texa[4] ),
    .B(\rbzero.texV[4] ),
    .Y(_03217_));
 sky130_fd_sc_hd__nand2_1 _20196_ (.A(\rbzero.traced_texa[4] ),
    .B(\rbzero.texV[4] ),
    .Y(_03218_));
 sky130_fd_sc_hd__and2b_1 _20197_ (.A_N(_03217_),
    .B(_03218_),
    .X(_03219_));
 sky130_fd_sc_hd__xnor2_1 _20198_ (.A(_03216_),
    .B(_03219_),
    .Y(_03220_));
 sky130_fd_sc_hd__a22o_1 _20199_ (.A1(\rbzero.texV[4] ),
    .A2(_03137_),
    .B1(_03142_),
    .B2(_03220_),
    .X(_01322_));
 sky130_fd_sc_hd__or2_1 _20200_ (.A(\rbzero.traced_texa[5] ),
    .B(\rbzero.texV[5] ),
    .X(_03221_));
 sky130_fd_sc_hd__nand2_1 _20201_ (.A(\rbzero.traced_texa[5] ),
    .B(\rbzero.texV[5] ),
    .Y(_03222_));
 sky130_fd_sc_hd__nand2_1 _20202_ (.A(_03221_),
    .B(_03222_),
    .Y(_03223_));
 sky130_fd_sc_hd__o21ai_1 _20203_ (.A1(_03216_),
    .A2(_03217_),
    .B1(_03218_),
    .Y(_03224_));
 sky130_fd_sc_hd__xnor2_1 _20204_ (.A(_03223_),
    .B(_03224_),
    .Y(_03225_));
 sky130_fd_sc_hd__a22o_1 _20205_ (.A1(\rbzero.texV[5] ),
    .A2(_03137_),
    .B1(_03142_),
    .B2(_03225_),
    .X(_01323_));
 sky130_fd_sc_hd__nor2_1 _20206_ (.A(\rbzero.traced_texa[6] ),
    .B(\rbzero.texV[6] ),
    .Y(_03226_));
 sky130_fd_sc_hd__nand2_1 _20207_ (.A(\rbzero.traced_texa[6] ),
    .B(\rbzero.texV[6] ),
    .Y(_03227_));
 sky130_fd_sc_hd__and2b_1 _20208_ (.A_N(_03226_),
    .B(_03227_),
    .X(_03228_));
 sky130_fd_sc_hd__a21boi_1 _20209_ (.A1(_03221_),
    .A2(_03224_),
    .B1_N(_03222_),
    .Y(_03229_));
 sky130_fd_sc_hd__xnor2_1 _20210_ (.A(_03228_),
    .B(_03229_),
    .Y(_03230_));
 sky130_fd_sc_hd__a22o_1 _20211_ (.A1(\rbzero.texV[6] ),
    .A2(_03137_),
    .B1(_03142_),
    .B2(_03230_),
    .X(_01324_));
 sky130_fd_sc_hd__xnor2_1 _20212_ (.A(\rbzero.traced_texa[7] ),
    .B(\rbzero.texV[7] ),
    .Y(_03231_));
 sky130_fd_sc_hd__o21ai_1 _20213_ (.A1(_03226_),
    .A2(_03229_),
    .B1(_03227_),
    .Y(_03232_));
 sky130_fd_sc_hd__xnor2_1 _20214_ (.A(_03231_),
    .B(_03232_),
    .Y(_03233_));
 sky130_fd_sc_hd__a22o_1 _20215_ (.A1(\rbzero.texV[7] ),
    .A2(_03137_),
    .B1(_03142_),
    .B2(_03233_),
    .X(_01325_));
 sky130_fd_sc_hd__nor2_1 _20216_ (.A(\rbzero.traced_texa[8] ),
    .B(\rbzero.texV[8] ),
    .Y(_03234_));
 sky130_fd_sc_hd__nand2_1 _20217_ (.A(\rbzero.traced_texa[8] ),
    .B(\rbzero.texV[8] ),
    .Y(_03235_));
 sky130_fd_sc_hd__and2b_1 _20218_ (.A_N(_03234_),
    .B(_03235_),
    .X(_03236_));
 sky130_fd_sc_hd__a21o_1 _20219_ (.A1(\rbzero.traced_texa[7] ),
    .A2(\rbzero.texV[7] ),
    .B1(_03232_),
    .X(_03237_));
 sky130_fd_sc_hd__o21ai_1 _20220_ (.A1(\rbzero.traced_texa[7] ),
    .A2(\rbzero.texV[7] ),
    .B1(_03237_),
    .Y(_03238_));
 sky130_fd_sc_hd__xnor2_1 _20221_ (.A(_03236_),
    .B(_03238_),
    .Y(_03239_));
 sky130_fd_sc_hd__a22o_1 _20222_ (.A1(\rbzero.texV[8] ),
    .A2(_03137_),
    .B1(_03142_),
    .B2(_03239_),
    .X(_01326_));
 sky130_fd_sc_hd__or2_1 _20223_ (.A(\rbzero.traced_texa[9] ),
    .B(\rbzero.texV[9] ),
    .X(_03240_));
 sky130_fd_sc_hd__nand2_1 _20224_ (.A(\rbzero.traced_texa[9] ),
    .B(\rbzero.texV[9] ),
    .Y(_03241_));
 sky130_fd_sc_hd__o21ai_1 _20225_ (.A1(_03234_),
    .A2(_03238_),
    .B1(_03235_),
    .Y(_03242_));
 sky130_fd_sc_hd__a21o_1 _20226_ (.A1(_03240_),
    .A2(_03241_),
    .B1(_03242_),
    .X(_03243_));
 sky130_fd_sc_hd__nand3_1 _20227_ (.A(_03240_),
    .B(_03241_),
    .C(_03242_),
    .Y(_03244_));
 sky130_fd_sc_hd__a32o_1 _20228_ (.A1(_09245_),
    .A2(_03243_),
    .A3(_03244_),
    .B1(_03064_),
    .B2(\rbzero.texV[9] ),
    .X(_01327_));
 sky130_fd_sc_hd__or2_1 _20229_ (.A(\rbzero.traced_texa[10] ),
    .B(\rbzero.texV[10] ),
    .X(_03245_));
 sky130_fd_sc_hd__nand2_1 _20230_ (.A(\rbzero.traced_texa[10] ),
    .B(\rbzero.texV[10] ),
    .Y(_03246_));
 sky130_fd_sc_hd__a21o_1 _20231_ (.A1(\rbzero.traced_texa[9] ),
    .A2(\rbzero.texV[9] ),
    .B1(_03242_),
    .X(_03247_));
 sky130_fd_sc_hd__a22o_1 _20232_ (.A1(_03245_),
    .A2(_03246_),
    .B1(_03247_),
    .B2(_03240_),
    .X(_03248_));
 sky130_fd_sc_hd__nand4_1 _20233_ (.A(_03240_),
    .B(_03245_),
    .C(_03246_),
    .D(_03247_),
    .Y(_03249_));
 sky130_fd_sc_hd__a32o_1 _20234_ (.A1(_09245_),
    .A2(_03248_),
    .A3(_03249_),
    .B1(_03064_),
    .B2(\rbzero.texV[10] ),
    .X(_01328_));
 sky130_fd_sc_hd__xnor2_1 _20235_ (.A(\rbzero.traced_texa[11] ),
    .B(\rbzero.texV[11] ),
    .Y(_03250_));
 sky130_fd_sc_hd__a21oi_1 _20236_ (.A1(_03246_),
    .A2(_03249_),
    .B1(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__a31o_1 _20237_ (.A1(_03246_),
    .A2(_03249_),
    .A3(_03250_),
    .B1(_09244_),
    .X(_03252_));
 sky130_fd_sc_hd__a2bb2o_1 _20238_ (.A1_N(_03251_),
    .A2_N(_03252_),
    .B1(\rbzero.texV[11] ),
    .B2(_03003_),
    .X(_01329_));
 sky130_fd_sc_hd__buf_4 _20239_ (.A(_03125_),
    .X(_03253_));
 sky130_fd_sc_hd__clkinv_2 _20240_ (.A(_03253_),
    .Y(_00337_));
 sky130_fd_sc_hd__clkinv_2 _20241_ (.A(_03253_),
    .Y(_00338_));
 sky130_fd_sc_hd__clkinv_2 _20242_ (.A(_03253_),
    .Y(_00339_));
 sky130_fd_sc_hd__clkinv_2 _20243_ (.A(_03253_),
    .Y(_00340_));
 sky130_fd_sc_hd__clkinv_2 _20244_ (.A(_03253_),
    .Y(_00341_));
 sky130_fd_sc_hd__clkinv_2 _20245_ (.A(_03253_),
    .Y(_00342_));
 sky130_fd_sc_hd__clkinv_2 _20246_ (.A(_03253_),
    .Y(_00343_));
 sky130_fd_sc_hd__clkinv_2 _20247_ (.A(_03253_),
    .Y(_00344_));
 sky130_fd_sc_hd__clkinv_2 _20248_ (.A(_03253_),
    .Y(_00345_));
 sky130_fd_sc_hd__clkinv_2 _20249_ (.A(_03253_),
    .Y(_00346_));
 sky130_fd_sc_hd__buf_4 _20250_ (.A(_03125_),
    .X(_03254_));
 sky130_fd_sc_hd__clkinv_2 _20251_ (.A(_03254_),
    .Y(_00347_));
 sky130_fd_sc_hd__clkinv_2 _20252_ (.A(_03254_),
    .Y(_00348_));
 sky130_fd_sc_hd__clkinv_2 _20253_ (.A(_03254_),
    .Y(_00349_));
 sky130_fd_sc_hd__clkinv_2 _20254_ (.A(_03254_),
    .Y(_00350_));
 sky130_fd_sc_hd__clkinv_2 _20255_ (.A(_03254_),
    .Y(_00351_));
 sky130_fd_sc_hd__clkinv_2 _20256_ (.A(_03254_),
    .Y(_00352_));
 sky130_fd_sc_hd__clkinv_2 _20257_ (.A(_03254_),
    .Y(_00353_));
 sky130_fd_sc_hd__clkinv_2 _20258_ (.A(_03254_),
    .Y(_00354_));
 sky130_fd_sc_hd__clkinv_2 _20259_ (.A(_03254_),
    .Y(_00355_));
 sky130_fd_sc_hd__clkinv_2 _20260_ (.A(_03254_),
    .Y(_00356_));
 sky130_fd_sc_hd__buf_4 _20261_ (.A(_03125_),
    .X(_03255_));
 sky130_fd_sc_hd__clkinv_2 _20262_ (.A(_03255_),
    .Y(_00357_));
 sky130_fd_sc_hd__clkinv_2 _20263_ (.A(_03255_),
    .Y(_00358_));
 sky130_fd_sc_hd__clkinv_2 _20264_ (.A(_03255_),
    .Y(_00359_));
 sky130_fd_sc_hd__clkinv_2 _20265_ (.A(_03255_),
    .Y(_00360_));
 sky130_fd_sc_hd__clkinv_2 _20266_ (.A(_03255_),
    .Y(_00361_));
 sky130_fd_sc_hd__clkinv_2 _20267_ (.A(_03255_),
    .Y(_00362_));
 sky130_fd_sc_hd__clkinv_2 _20268_ (.A(_03255_),
    .Y(_00363_));
 sky130_fd_sc_hd__clkinv_2 _20269_ (.A(_03255_),
    .Y(_00364_));
 sky130_fd_sc_hd__clkinv_2 _20270_ (.A(_03255_),
    .Y(_00365_));
 sky130_fd_sc_hd__clkinv_2 _20271_ (.A(_03255_),
    .Y(_00366_));
 sky130_fd_sc_hd__buf_4 _20272_ (.A(_03125_),
    .X(_03256_));
 sky130_fd_sc_hd__clkinv_2 _20273_ (.A(_03256_),
    .Y(_00367_));
 sky130_fd_sc_hd__clkinv_2 _20274_ (.A(_03256_),
    .Y(_00368_));
 sky130_fd_sc_hd__clkinv_2 _20275_ (.A(_03256_),
    .Y(_00369_));
 sky130_fd_sc_hd__clkinv_2 _20276_ (.A(_03256_),
    .Y(_00370_));
 sky130_fd_sc_hd__clkinv_2 _20277_ (.A(_03256_),
    .Y(_00371_));
 sky130_fd_sc_hd__clkinv_2 _20278_ (.A(_03256_),
    .Y(_00372_));
 sky130_fd_sc_hd__clkinv_2 _20279_ (.A(_03256_),
    .Y(_00373_));
 sky130_fd_sc_hd__clkinv_2 _20280_ (.A(_03256_),
    .Y(_00374_));
 sky130_fd_sc_hd__clkinv_2 _20281_ (.A(_03256_),
    .Y(_00375_));
 sky130_fd_sc_hd__clkinv_2 _20282_ (.A(_03256_),
    .Y(_00376_));
 sky130_fd_sc_hd__buf_4 _20283_ (.A(_04702_),
    .X(_03257_));
 sky130_fd_sc_hd__clkinv_2 _20284_ (.A(_03257_),
    .Y(_00377_));
 sky130_fd_sc_hd__clkinv_2 _20285_ (.A(_03257_),
    .Y(_00378_));
 sky130_fd_sc_hd__clkinv_2 _20286_ (.A(_03257_),
    .Y(_00379_));
 sky130_fd_sc_hd__clkinv_2 _20287_ (.A(_03257_),
    .Y(_00380_));
 sky130_fd_sc_hd__clkinv_2 _20288_ (.A(_03257_),
    .Y(_00381_));
 sky130_fd_sc_hd__clkinv_2 _20289_ (.A(_03257_),
    .Y(_00382_));
 sky130_fd_sc_hd__clkinv_2 _20290_ (.A(_03257_),
    .Y(_00383_));
 sky130_fd_sc_hd__clkinv_2 _20291_ (.A(_03257_),
    .Y(_00384_));
 sky130_fd_sc_hd__clkinv_2 _20292_ (.A(_03257_),
    .Y(_00385_));
 sky130_fd_sc_hd__clkinv_2 _20293_ (.A(_03257_),
    .Y(_00386_));
 sky130_fd_sc_hd__buf_4 _20294_ (.A(_04702_),
    .X(_03258_));
 sky130_fd_sc_hd__clkinv_2 _20295_ (.A(_03258_),
    .Y(_00387_));
 sky130_fd_sc_hd__clkinv_2 _20296_ (.A(_03258_),
    .Y(_00388_));
 sky130_fd_sc_hd__clkinv_2 _20297_ (.A(_03258_),
    .Y(_00389_));
 sky130_fd_sc_hd__clkinv_2 _20298_ (.A(_03258_),
    .Y(_00390_));
 sky130_fd_sc_hd__clkinv_2 _20299_ (.A(_03258_),
    .Y(_00391_));
 sky130_fd_sc_hd__clkinv_2 _20300_ (.A(_03258_),
    .Y(_00392_));
 sky130_fd_sc_hd__clkinv_2 _20301_ (.A(_03258_),
    .Y(_00393_));
 sky130_fd_sc_hd__clkinv_2 _20302_ (.A(_03258_),
    .Y(_00394_));
 sky130_fd_sc_hd__clkinv_2 _20303_ (.A(_03258_),
    .Y(_00395_));
 sky130_fd_sc_hd__clkinv_2 _20304_ (.A(_03258_),
    .Y(_00396_));
 sky130_fd_sc_hd__clkinv_2 _20305_ (.A(_02855_),
    .Y(_00397_));
 sky130_fd_sc_hd__clkinv_2 _20306_ (.A(_02855_),
    .Y(_00398_));
 sky130_fd_sc_hd__clkinv_2 _20307_ (.A(_02855_),
    .Y(_00399_));
 sky130_fd_sc_hd__clkinv_2 _20308_ (.A(_02855_),
    .Y(_00400_));
 sky130_fd_sc_hd__o2bb2ai_1 _20309_ (.A1_N(\rbzero.traced_texVinit[0] ),
    .A2_N(_09255_),
    .B1(_08573_),
    .B2(_09269_),
    .Y(_01394_));
 sky130_fd_sc_hd__a22o_1 _20310_ (.A1(\rbzero.traced_texVinit[1] ),
    .A2(_09266_),
    .B1(_08571_),
    .B2(_09261_),
    .X(_01395_));
 sky130_fd_sc_hd__a22o_1 _20311_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(_09266_),
    .B1(_08564_),
    .B2(_09261_),
    .X(_01396_));
 sky130_fd_sc_hd__a2bb2o_1 _20312_ (.A1_N(_08700_),
    .A2_N(_09269_),
    .B1(\rbzero.traced_texVinit[3] ),
    .B2(_09255_),
    .X(_01397_));
 sky130_fd_sc_hd__inv_2 _20313_ (.A(_08828_),
    .Y(_03259_));
 sky130_fd_sc_hd__a22o_1 _20314_ (.A1(\rbzero.traced_texVinit[4] ),
    .A2(_09266_),
    .B1(_03259_),
    .B2(_09261_),
    .X(_01398_));
 sky130_fd_sc_hd__a22o_1 _20315_ (.A1(\rbzero.traced_texVinit[5] ),
    .A2(_09266_),
    .B1(_08959_),
    .B2(_09261_),
    .X(_01399_));
 sky130_fd_sc_hd__a22o_1 _20316_ (.A1(\rbzero.traced_texVinit[6] ),
    .A2(_09266_),
    .B1(_09099_),
    .B2(_09261_),
    .X(_01400_));
 sky130_fd_sc_hd__a22o_1 _20317_ (.A1(\rbzero.traced_texVinit[7] ),
    .A2(_09266_),
    .B1(_09237_),
    .B2(_09261_),
    .X(_01401_));
 sky130_fd_sc_hd__clkbuf_4 _20318_ (.A(_02197_),
    .X(_03260_));
 sky130_fd_sc_hd__a22o_1 _20319_ (.A1(\rbzero.traced_texVinit[8] ),
    .A2(_03260_),
    .B1(_09267_),
    .B2(_09507_),
    .X(_01402_));
 sky130_fd_sc_hd__a22o_1 _20320_ (.A1(\rbzero.traced_texVinit[9] ),
    .A2(_03260_),
    .B1(_09267_),
    .B2(_09640_),
    .X(_01403_));
 sky130_fd_sc_hd__a22o_1 _20321_ (.A1(\rbzero.traced_texVinit[10] ),
    .A2(_03260_),
    .B1(_09267_),
    .B2(_09764_),
    .X(_01404_));
 sky130_fd_sc_hd__a22o_1 _20322_ (.A1(\rbzero.traced_texVinit[11] ),
    .A2(_03260_),
    .B1(_09267_),
    .B2(_09887_),
    .X(_01405_));
 sky130_fd_sc_hd__nor2_1 _20323_ (.A(\gpout0.clk_div[0] ),
    .B(_03003_),
    .Y(_01406_));
 sky130_fd_sc_hd__nand2_1 _20324_ (.A(\gpout0.clk_div[0] ),
    .B(\gpout0.clk_div[1] ),
    .Y(_03261_));
 sky130_fd_sc_hd__or2_1 _20325_ (.A(\gpout0.clk_div[0] ),
    .B(\gpout0.clk_div[1] ),
    .X(_03262_));
 sky130_fd_sc_hd__and3_1 _20326_ (.A(_09247_),
    .B(_03261_),
    .C(_03262_),
    .X(_03263_));
 sky130_fd_sc_hd__clkbuf_1 _20327_ (.A(_03263_),
    .X(_01407_));
 sky130_fd_sc_hd__nor2_1 _20328_ (.A(\gpout1.clk_div[0] ),
    .B(_03003_),
    .Y(_01408_));
 sky130_fd_sc_hd__nand2_1 _20329_ (.A(\gpout1.clk_div[0] ),
    .B(\gpout1.clk_div[1] ),
    .Y(_03264_));
 sky130_fd_sc_hd__or2_1 _20330_ (.A(\gpout1.clk_div[0] ),
    .B(\gpout1.clk_div[1] ),
    .X(_03265_));
 sky130_fd_sc_hd__and3_1 _20331_ (.A(_02727_),
    .B(_03264_),
    .C(_03265_),
    .X(_03266_));
 sky130_fd_sc_hd__clkbuf_1 _20332_ (.A(_03266_),
    .X(_01409_));
 sky130_fd_sc_hd__or2_1 _20333_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-9] ),
    .X(_03267_));
 sky130_fd_sc_hd__a32o_1 _20334_ (.A1(_02287_),
    .A2(_02148_),
    .A3(_03267_),
    .B1(_03260_),
    .B2(\rbzero.wall_tracer.rayAddendX[-9] ),
    .X(_01410_));
 sky130_fd_sc_hd__a21bo_1 _20335_ (.A1(_02147_),
    .A2(_02149_),
    .B1_N(_02148_),
    .X(_03268_));
 sky130_fd_sc_hd__a32o_1 _20336_ (.A1(_02287_),
    .A2(_02150_),
    .A3(_03268_),
    .B1(_03260_),
    .B2(\rbzero.wall_tracer.rayAddendX[-8] ),
    .X(_01411_));
 sky130_fd_sc_hd__and2b_1 _20337_ (.A_N(_02146_),
    .B(_02152_),
    .X(_03269_));
 sky130_fd_sc_hd__xnor2_1 _20338_ (.A(_02151_),
    .B(_03269_),
    .Y(_03270_));
 sky130_fd_sc_hd__a22o_1 _20339_ (.A1(\rbzero.wall_tracer.rayAddendX[-7] ),
    .A2(_03260_),
    .B1(_09267_),
    .B2(_03270_),
    .X(_01412_));
 sky130_fd_sc_hd__xnor2_1 _20340_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[-6] ),
    .Y(_03271_));
 sky130_fd_sc_hd__xnor2_1 _20341_ (.A(_02153_),
    .B(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__a22o_1 _20342_ (.A1(\rbzero.wall_tracer.rayAddendX[-6] ),
    .A2(_03260_),
    .B1(_09267_),
    .B2(_03272_),
    .X(_01413_));
 sky130_fd_sc_hd__or2_1 _20343_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-9] ),
    .X(_03273_));
 sky130_fd_sc_hd__a32o_1 _20344_ (.A1(_09257_),
    .A2(_02375_),
    .A3(_03273_),
    .B1(_02158_),
    .B2(\rbzero.wall_tracer.rayAddendY[-9] ),
    .X(_01414_));
 sky130_fd_sc_hd__a21bo_1 _20345_ (.A1(_02374_),
    .A2(_02376_),
    .B1_N(_02375_),
    .X(_03274_));
 sky130_fd_sc_hd__a32o_1 _20346_ (.A1(_09257_),
    .A2(_02377_),
    .A3(_03274_),
    .B1(_02158_),
    .B2(\rbzero.wall_tracer.rayAddendY[-8] ),
    .X(_01415_));
 sky130_fd_sc_hd__and2b_1 _20347_ (.A_N(_02373_),
    .B(_02379_),
    .X(_03275_));
 sky130_fd_sc_hd__xnor2_1 _20348_ (.A(_02378_),
    .B(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__a22o_1 _20349_ (.A1(\rbzero.wall_tracer.rayAddendY[-7] ),
    .A2(_03260_),
    .B1(_09267_),
    .B2(_03276_),
    .X(_01416_));
 sky130_fd_sc_hd__xnor2_1 _20350_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[-6] ),
    .Y(_03277_));
 sky130_fd_sc_hd__xnor2_1 _20351_ (.A(_02380_),
    .B(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__a22o_1 _20352_ (.A1(\rbzero.wall_tracer.rayAddendY[-6] ),
    .A2(_03260_),
    .B1(_09267_),
    .B2(_03278_),
    .X(_01417_));
 sky130_fd_sc_hd__nor2_1 _20353_ (.A(\gpout2.clk_div[0] ),
    .B(_03003_),
    .Y(_01418_));
 sky130_fd_sc_hd__nand2_1 _20354_ (.A(\gpout2.clk_div[0] ),
    .B(\gpout2.clk_div[1] ),
    .Y(_03279_));
 sky130_fd_sc_hd__or2_1 _20355_ (.A(\gpout2.clk_div[0] ),
    .B(\gpout2.clk_div[1] ),
    .X(_03280_));
 sky130_fd_sc_hd__and3_1 _20356_ (.A(_02727_),
    .B(_03279_),
    .C(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__clkbuf_1 _20357_ (.A(_03281_),
    .X(_01419_));
 sky130_fd_sc_hd__nor2_1 _20358_ (.A(\gpout3.clk_div[0] ),
    .B(_03003_),
    .Y(_01420_));
 sky130_fd_sc_hd__nand2_1 _20359_ (.A(\gpout3.clk_div[1] ),
    .B(\gpout3.clk_div[0] ),
    .Y(_03282_));
 sky130_fd_sc_hd__or2_1 _20360_ (.A(\gpout3.clk_div[1] ),
    .B(\gpout3.clk_div[0] ),
    .X(_03283_));
 sky130_fd_sc_hd__and3_1 _20361_ (.A(_02727_),
    .B(_03282_),
    .C(_03283_),
    .X(_03284_));
 sky130_fd_sc_hd__clkbuf_1 _20362_ (.A(_03284_),
    .X(_01421_));
 sky130_fd_sc_hd__nor2_1 _20363_ (.A(\gpout4.clk_div[0] ),
    .B(_03003_),
    .Y(_01422_));
 sky130_fd_sc_hd__nand2_1 _20364_ (.A(\gpout4.clk_div[1] ),
    .B(\gpout4.clk_div[0] ),
    .Y(_03285_));
 sky130_fd_sc_hd__or2_1 _20365_ (.A(\gpout4.clk_div[1] ),
    .B(\gpout4.clk_div[0] ),
    .X(_03286_));
 sky130_fd_sc_hd__and3_1 _20366_ (.A(_02727_),
    .B(_03285_),
    .C(_03286_),
    .X(_03287_));
 sky130_fd_sc_hd__clkbuf_1 _20367_ (.A(_03287_),
    .X(_01423_));
 sky130_fd_sc_hd__dfxtp_2 _20368_ (.CLK(net92),
    .D(_00401_),
    .Q(\rbzero.map_rom.d6 ));
 sky130_fd_sc_hd__dfxtp_2 _20369_ (.CLK(net92),
    .D(_00402_),
    .Q(\rbzero.map_rom.c6 ));
 sky130_fd_sc_hd__dfxtp_1 _20370_ (.CLK(net97),
    .D(_00403_),
    .Q(\rbzero.map_rom.b6 ));
 sky130_fd_sc_hd__dfxtp_2 _20371_ (.CLK(net92),
    .D(_00404_),
    .Q(\rbzero.map_rom.a6 ));
 sky130_fd_sc_hd__dfxtp_1 _20372_ (.CLK(net97),
    .D(_00405_),
    .Q(\rbzero.map_rom.i_row[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20373_ (.CLK(net118),
    .D(_00011_),
    .Q(\rbzero.wall_tracer.rcp_sel[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20374_ (.CLK(net118),
    .D(_00012_),
    .Q(\rbzero.wall_tracer.rcp_sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20375_ (.CLK(net126),
    .D(_00406_),
    .Q(\rbzero.wall_tracer.stepDistY[-12] ));
 sky130_fd_sc_hd__dfxtp_1 _20376_ (.CLK(net124),
    .D(_00407_),
    .Q(\rbzero.wall_tracer.stepDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20377_ (.CLK(net120),
    .D(_00408_),
    .Q(\rbzero.wall_tracer.stepDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20378_ (.CLK(net116),
    .D(_00409_),
    .Q(\rbzero.wall_tracer.stepDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20379_ (.CLK(net116),
    .D(_00410_),
    .Q(\rbzero.wall_tracer.stepDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20380_ (.CLK(net116),
    .D(_00411_),
    .Q(\rbzero.wall_tracer.stepDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20381_ (.CLK(net116),
    .D(_00412_),
    .Q(\rbzero.wall_tracer.stepDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20382_ (.CLK(net121),
    .D(_00413_),
    .Q(\rbzero.wall_tracer.stepDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20383_ (.CLK(net121),
    .D(_00414_),
    .Q(\rbzero.wall_tracer.stepDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20384_ (.CLK(net131),
    .D(_00415_),
    .Q(\rbzero.wall_tracer.stepDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20385_ (.CLK(net131),
    .D(_00416_),
    .Q(\rbzero.wall_tracer.stepDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20386_ (.CLK(net131),
    .D(_00417_),
    .Q(\rbzero.wall_tracer.stepDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20387_ (.CLK(net135),
    .D(_00418_),
    .Q(\rbzero.wall_tracer.stepDistY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20388_ (.CLK(net135),
    .D(_00419_),
    .Q(\rbzero.wall_tracer.stepDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20389_ (.CLK(net135),
    .D(_00420_),
    .Q(\rbzero.wall_tracer.stepDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20390_ (.CLK(net135),
    .D(_00421_),
    .Q(\rbzero.wall_tracer.stepDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20391_ (.CLK(net135),
    .D(_00422_),
    .Q(\rbzero.wall_tracer.stepDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20392_ (.CLK(net138),
    .D(_00423_),
    .Q(\rbzero.wall_tracer.stepDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20393_ (.CLK(net138),
    .D(_00424_),
    .Q(\rbzero.wall_tracer.stepDistY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20394_ (.CLK(net138),
    .D(_00425_),
    .Q(\rbzero.wall_tracer.stepDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20395_ (.CLK(net137),
    .D(_00426_),
    .Q(\rbzero.wall_tracer.stepDistY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20396_ (.CLK(net138),
    .D(_00427_),
    .Q(\rbzero.wall_tracer.stepDistY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20397_ (.CLK(net138),
    .D(_00428_),
    .Q(\rbzero.wall_tracer.stepDistY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20398_ (.CLK(net125),
    .D(_00429_),
    .Q(\rbzero.wall_tracer.stepDistY[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20399_ (.CLK(net121),
    .D(_00430_),
    .Q(\rbzero.wall_tracer.visualWallDist[-12] ));
 sky130_fd_sc_hd__dfxtp_2 _20400_ (.CLK(net123),
    .D(_00431_),
    .Q(\rbzero.wall_tracer.visualWallDist[-11] ));
 sky130_fd_sc_hd__dfxtp_4 _20401_ (.CLK(net121),
    .D(_00432_),
    .Q(\rbzero.wall_tracer.visualWallDist[-10] ));
 sky130_fd_sc_hd__dfxtp_2 _20402_ (.CLK(net121),
    .D(_00433_),
    .Q(\rbzero.wall_tracer.visualWallDist[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _20403_ (.CLK(net121),
    .D(_00434_),
    .Q(\rbzero.wall_tracer.visualWallDist[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _20404_ (.CLK(net119),
    .D(_00435_),
    .Q(\rbzero.wall_tracer.visualWallDist[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _20405_ (.CLK(net119),
    .D(_00436_),
    .Q(\rbzero.wall_tracer.visualWallDist[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _20406_ (.CLK(net128),
    .D(_00437_),
    .Q(\rbzero.wall_tracer.visualWallDist[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _20407_ (.CLK(net128),
    .D(_00438_),
    .Q(\rbzero.wall_tracer.visualWallDist[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20408_ (.CLK(net130),
    .D(_00439_),
    .Q(\rbzero.wall_tracer.visualWallDist[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _20409_ (.CLK(net130),
    .D(_00440_),
    .Q(\rbzero.wall_tracer.visualWallDist[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _20410_ (.CLK(net130),
    .D(_00441_),
    .Q(\rbzero.wall_tracer.visualWallDist[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _20411_ (.CLK(net130),
    .D(_00442_),
    .Q(\rbzero.wall_tracer.visualWallDist[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20412_ (.CLK(net130),
    .D(_00443_),
    .Q(\rbzero.wall_tracer.visualWallDist[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20413_ (.CLK(net130),
    .D(_00444_),
    .Q(\rbzero.wall_tracer.visualWallDist[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20414_ (.CLK(net136),
    .D(_00445_),
    .Q(\rbzero.wall_tracer.visualWallDist[3] ));
 sky130_fd_sc_hd__dfxtp_4 _20415_ (.CLK(net136),
    .D(_00446_),
    .Q(\rbzero.wall_tracer.visualWallDist[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20416_ (.CLK(net135),
    .D(_00447_),
    .Q(\rbzero.wall_tracer.visualWallDist[5] ));
 sky130_fd_sc_hd__dfxtp_4 _20417_ (.CLK(net136),
    .D(_00448_),
    .Q(\rbzero.wall_tracer.visualWallDist[6] ));
 sky130_fd_sc_hd__dfxtp_4 _20418_ (.CLK(net136),
    .D(_00449_),
    .Q(\rbzero.wall_tracer.visualWallDist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20419_ (.CLK(net128),
    .D(_00450_),
    .Q(\rbzero.wall_tracer.visualWallDist[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20420_ (.CLK(net123),
    .D(_00451_),
    .Q(\rbzero.wall_tracer.visualWallDist[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20421_ (.CLK(net130),
    .D(_00452_),
    .Q(\rbzero.wall_tracer.visualWallDist[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20422_ (.CLK(net123),
    .D(_00453_),
    .Q(\rbzero.wall_tracer.visualWallDist[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20423_ (.CLK(net126),
    .D(_00454_),
    .Q(\rbzero.wall_tracer.stepDistX[-12] ));
 sky130_fd_sc_hd__dfxtp_1 _20424_ (.CLK(net124),
    .D(_00455_),
    .Q(\rbzero.wall_tracer.stepDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20425_ (.CLK(net117),
    .D(_00456_),
    .Q(\rbzero.wall_tracer.stepDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20426_ (.CLK(net117),
    .D(_00457_),
    .Q(\rbzero.wall_tracer.stepDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20427_ (.CLK(net117),
    .D(_00458_),
    .Q(\rbzero.wall_tracer.stepDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20428_ (.CLK(net118),
    .D(_00459_),
    .Q(\rbzero.wall_tracer.stepDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20429_ (.CLK(net117),
    .D(_00460_),
    .Q(\rbzero.wall_tracer.stepDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20430_ (.CLK(net119),
    .D(_00461_),
    .Q(\rbzero.wall_tracer.stepDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20431_ (.CLK(net121),
    .D(_00462_),
    .Q(\rbzero.wall_tracer.stepDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20432_ (.CLK(net131),
    .D(_00463_),
    .Q(\rbzero.wall_tracer.stepDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20433_ (.CLK(net131),
    .D(_00464_),
    .Q(\rbzero.wall_tracer.stepDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20434_ (.CLK(net131),
    .D(_00465_),
    .Q(\rbzero.wall_tracer.stepDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _20435_ (.CLK(net135),
    .D(_00466_),
    .Q(\rbzero.wall_tracer.stepDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20436_ (.CLK(net135),
    .D(_00467_),
    .Q(\rbzero.wall_tracer.stepDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20437_ (.CLK(net135),
    .D(_00468_),
    .Q(\rbzero.wall_tracer.stepDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20438_ (.CLK(net139),
    .D(_00469_),
    .Q(\rbzero.wall_tracer.stepDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20439_ (.CLK(net138),
    .D(_00470_),
    .Q(\rbzero.wall_tracer.stepDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20440_ (.CLK(net138),
    .D(_00471_),
    .Q(\rbzero.wall_tracer.stepDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20441_ (.CLK(net138),
    .D(_00472_),
    .Q(\rbzero.wall_tracer.stepDistX[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20442_ (.CLK(net138),
    .D(_00473_),
    .Q(\rbzero.wall_tracer.stepDistX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20443_ (.CLK(net137),
    .D(_00474_),
    .Q(\rbzero.wall_tracer.stepDistX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20444_ (.CLK(net138),
    .D(_00475_),
    .Q(\rbzero.wall_tracer.stepDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20445_ (.CLK(net139),
    .D(_00476_),
    .Q(\rbzero.wall_tracer.stepDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20446_ (.CLK(net125),
    .D(_00477_),
    .Q(\rbzero.wall_tracer.stepDistX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20447_ (.CLK(net95),
    .D(_00013_),
    .Q(\rbzero.wall_tracer.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20448_ (.CLK(net123),
    .D(_00015_),
    .Q(\rbzero.wall_tracer.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20449_ (.CLK(net118),
    .D(_00000_),
    .Q(\rbzero.wall_tracer.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20450_ (.CLK(net118),
    .D(_00001_),
    .Q(\rbzero.wall_tracer.state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20451_ (.CLK(net119),
    .D(_00002_),
    .Q(\rbzero.wall_tracer.state[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20452_ (.CLK(net118),
    .D(_00003_),
    .Q(\rbzero.wall_tracer.state[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20453_ (.CLK(net117),
    .D(_00004_),
    .Q(\rbzero.wall_tracer.state[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20454_ (.CLK(net118),
    .D(_00005_),
    .Q(\rbzero.wall_tracer.state[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20455_ (.CLK(net97),
    .D(_00016_),
    .Q(\rbzero.wall_tracer.state[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20456_ (.CLK(net119),
    .D(_00006_),
    .Q(\rbzero.wall_tracer.state[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20457_ (.CLK(net94),
    .D(_00007_),
    .Q(\rbzero.wall_tracer.state[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20458_ (.CLK(net118),
    .D(_00008_),
    .Q(\rbzero.wall_tracer.state[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20459_ (.CLK(net118),
    .D(_00009_),
    .Q(\rbzero.wall_tracer.state[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20460_ (.CLK(net126),
    .D(_00010_),
    .Q(\rbzero.wall_tracer.state[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20461_ (.CLK(net94),
    .D(_00014_),
    .Q(\rbzero.wall_tracer.state[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20462_ (.CLK(net96),
    .D(_00478_),
    .Q(\rbzero.wall_tracer.wall[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20463_ (.CLK(net96),
    .D(_00479_),
    .Q(\rbzero.wall_tracer.wall[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20464_ (.CLK(net118),
    .D(_00480_),
    .Q(\rbzero.wall_tracer.side ));
 sky130_fd_sc_hd__dfxtp_1 _20465_ (.CLK(net128),
    .D(_00481_),
    .Q(\rbzero.wall_tracer.texu[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20466_ (.CLK(net119),
    .D(_00482_),
    .Q(\rbzero.wall_tracer.texu[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20467_ (.CLK(net127),
    .D(_00483_),
    .Q(\rbzero.wall_tracer.texu[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20468_ (.CLK(net119),
    .D(_00484_),
    .Q(\rbzero.wall_tracer.texu[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20469_ (.CLK(net119),
    .D(_00485_),
    .Q(\rbzero.wall_tracer.texu[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20470_ (.CLK(net119),
    .D(_00486_),
    .Q(\rbzero.wall_tracer.texu[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20471_ (.CLK(net111),
    .D(_00487_),
    .Q(\gpout0.hpos[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20472_ (.CLK(net111),
    .D(_00488_),
    .Q(\gpout0.hpos[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20473_ (.CLK(net112),
    .D(_00489_),
    .Q(\gpout0.hpos[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20474_ (.CLK(net94),
    .D(_00490_),
    .Q(\gpout0.hpos[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20475_ (.CLK(net96),
    .D(_00491_),
    .Q(\gpout0.hpos[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20476_ (.CLK(net96),
    .D(_00492_),
    .Q(\gpout0.hpos[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20477_ (.CLK(net96),
    .D(_00493_),
    .Q(\gpout0.hpos[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20478_ (.CLK(net94),
    .D(_00494_),
    .Q(\gpout0.hpos[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20479_ (.CLK(net94),
    .D(_00495_),
    .Q(\gpout0.hpos[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20480_ (.CLK(net94),
    .D(_00496_),
    .Q(\gpout0.hpos[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20481_ (.CLK(net96),
    .D(_00497_),
    .Q(\rbzero.row_render.side ));
 sky130_fd_sc_hd__dfxtp_1 _20482_ (.CLK(net111),
    .D(_00498_),
    .Q(\rbzero.row_render.size[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20483_ (.CLK(net111),
    .D(_00499_),
    .Q(\rbzero.row_render.size[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20484_ (.CLK(net111),
    .D(_00500_),
    .Q(\rbzero.row_render.size[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20485_ (.CLK(net111),
    .D(_00501_),
    .Q(\rbzero.row_render.size[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20486_ (.CLK(net112),
    .D(_00502_),
    .Q(\rbzero.row_render.size[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20487_ (.CLK(net112),
    .D(_00503_),
    .Q(\rbzero.row_render.size[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20488_ (.CLK(net112),
    .D(_00504_),
    .Q(\rbzero.row_render.size[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20489_ (.CLK(net112),
    .D(_00505_),
    .Q(\rbzero.row_render.size[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20490_ (.CLK(net112),
    .D(_00506_),
    .Q(\rbzero.row_render.size[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20491_ (.CLK(net114),
    .D(_00507_),
    .Q(\rbzero.row_render.size[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20492_ (.CLK(net114),
    .D(_00508_),
    .Q(\rbzero.row_render.size[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20493_ (.CLK(net111),
    .D(_00509_),
    .Q(\rbzero.row_render.texu[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20494_ (.CLK(net111),
    .D(_00510_),
    .Q(\rbzero.row_render.texu[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20495_ (.CLK(net127),
    .D(_00511_),
    .Q(\rbzero.row_render.texu[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20496_ (.CLK(net127),
    .D(_00512_),
    .Q(\rbzero.row_render.texu[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20497_ (.CLK(net127),
    .D(_00513_),
    .Q(\rbzero.row_render.texu[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20498_ (.CLK(net127),
    .D(_00514_),
    .Q(\rbzero.row_render.texu[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20499_ (.CLK(net128),
    .D(_00515_),
    .Q(\rbzero.traced_texa[-12] ));
 sky130_fd_sc_hd__dfxtp_1 _20500_ (.CLK(net128),
    .D(_00516_),
    .Q(\rbzero.traced_texa[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20501_ (.CLK(net133),
    .D(_00517_),
    .Q(\rbzero.traced_texa[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20502_ (.CLK(net129),
    .D(_00518_),
    .Q(\rbzero.traced_texa[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20503_ (.CLK(net133),
    .D(_00519_),
    .Q(\rbzero.traced_texa[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20504_ (.CLK(net132),
    .D(_00520_),
    .Q(\rbzero.traced_texa[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20505_ (.CLK(net133),
    .D(_00521_),
    .Q(\rbzero.traced_texa[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20506_ (.CLK(net132),
    .D(_00522_),
    .Q(\rbzero.traced_texa[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20507_ (.CLK(net132),
    .D(_00523_),
    .Q(\rbzero.traced_texa[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20508_ (.CLK(net132),
    .D(_00524_),
    .Q(\rbzero.traced_texa[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20509_ (.CLK(net129),
    .D(_00525_),
    .Q(\rbzero.traced_texa[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20510_ (.CLK(net132),
    .D(_00526_),
    .Q(\rbzero.traced_texa[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20511_ (.CLK(net128),
    .D(_00527_),
    .Q(\rbzero.traced_texa[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20512_ (.CLK(net127),
    .D(_00528_),
    .Q(\rbzero.traced_texa[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20513_ (.CLK(net127),
    .D(_00529_),
    .Q(\rbzero.traced_texa[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20514_ (.CLK(net129),
    .D(_00530_),
    .Q(\rbzero.traced_texa[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20515_ (.CLK(net129),
    .D(_00531_),
    .Q(\rbzero.traced_texa[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20516_ (.CLK(net132),
    .D(_00532_),
    .Q(\rbzero.traced_texa[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20517_ (.CLK(net132),
    .D(_00533_),
    .Q(\rbzero.traced_texa[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20518_ (.CLK(net132),
    .D(_00534_),
    .Q(\rbzero.traced_texa[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20519_ (.CLK(net129),
    .D(_00535_),
    .Q(\rbzero.traced_texa[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20520_ (.CLK(net129),
    .D(_00536_),
    .Q(\rbzero.traced_texa[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20521_ (.CLK(net113),
    .D(_00537_),
    .Q(\rbzero.traced_texa[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20522_ (.CLK(net113),
    .D(_00538_),
    .Q(\rbzero.traced_texa[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20523_ (.CLK(net96),
    .D(_00539_),
    .Q(\rbzero.row_render.wall[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20524_ (.CLK(net96),
    .D(_00540_),
    .Q(\rbzero.row_render.wall[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20525_ (.CLK(net124),
    .D(_00541_),
    .Q(\rbzero.wall_tracer.trackDistX[-12] ));
 sky130_fd_sc_hd__dfxtp_1 _20526_ (.CLK(net123),
    .D(_00542_),
    .Q(\rbzero.wall_tracer.trackDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20527_ (.CLK(net120),
    .D(_00543_),
    .Q(\rbzero.wall_tracer.trackDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20528_ (.CLK(net120),
    .D(_00544_),
    .Q(\rbzero.wall_tracer.trackDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20529_ (.CLK(net120),
    .D(_00545_),
    .Q(\rbzero.wall_tracer.trackDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20530_ (.CLK(net120),
    .D(_00546_),
    .Q(\rbzero.wall_tracer.trackDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20531_ (.CLK(net121),
    .D(_00547_),
    .Q(\rbzero.wall_tracer.trackDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20532_ (.CLK(net121),
    .D(_00548_),
    .Q(\rbzero.wall_tracer.trackDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20533_ (.CLK(net123),
    .D(_00549_),
    .Q(\rbzero.wall_tracer.trackDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20534_ (.CLK(net130),
    .D(_00550_),
    .Q(\rbzero.wall_tracer.trackDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20535_ (.CLK(net131),
    .D(_00551_),
    .Q(\rbzero.wall_tracer.trackDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20536_ (.CLK(net131),
    .D(_00552_),
    .Q(\rbzero.wall_tracer.trackDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20537_ (.CLK(net136),
    .D(_00553_),
    .Q(\rbzero.wall_tracer.trackDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20538_ (.CLK(net135),
    .D(_00554_),
    .Q(\rbzero.wall_tracer.trackDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20539_ (.CLK(net139),
    .D(_00555_),
    .Q(\rbzero.wall_tracer.trackDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20540_ (.CLK(net123),
    .D(_00556_),
    .Q(\rbzero.wall_tracer.trackDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20541_ (.CLK(net137),
    .D(_00557_),
    .Q(\rbzero.wall_tracer.trackDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20542_ (.CLK(net137),
    .D(_00558_),
    .Q(\rbzero.wall_tracer.trackDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20543_ (.CLK(net137),
    .D(_00559_),
    .Q(\rbzero.wall_tracer.trackDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20544_ (.CLK(net137),
    .D(_00560_),
    .Q(\rbzero.wall_tracer.trackDistX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20545_ (.CLK(net137),
    .D(_00561_),
    .Q(\rbzero.wall_tracer.trackDistX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20546_ (.CLK(net125),
    .D(_00562_),
    .Q(\rbzero.wall_tracer.trackDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20547_ (.CLK(net125),
    .D(_00563_),
    .Q(\rbzero.wall_tracer.trackDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20548_ (.CLK(net123),
    .D(_00564_),
    .Q(\rbzero.wall_tracer.trackDistX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20549_ (.CLK(net124),
    .D(_00565_),
    .Q(\rbzero.wall_tracer.trackDistY[-12] ));
 sky130_fd_sc_hd__dfxtp_1 _20550_ (.CLK(net124),
    .D(_00566_),
    .Q(\rbzero.wall_tracer.trackDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20551_ (.CLK(net120),
    .D(_00567_),
    .Q(\rbzero.wall_tracer.trackDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20552_ (.CLK(net120),
    .D(_00568_),
    .Q(\rbzero.wall_tracer.trackDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20553_ (.CLK(net120),
    .D(_00569_),
    .Q(\rbzero.wall_tracer.trackDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20554_ (.CLK(net120),
    .D(_00570_),
    .Q(\rbzero.wall_tracer.trackDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20555_ (.CLK(net120),
    .D(_00571_),
    .Q(\rbzero.wall_tracer.trackDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20556_ (.CLK(net121),
    .D(_00572_),
    .Q(\rbzero.wall_tracer.trackDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20557_ (.CLK(net123),
    .D(_00573_),
    .Q(\rbzero.wall_tracer.trackDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20558_ (.CLK(net136),
    .D(_00574_),
    .Q(\rbzero.wall_tracer.trackDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20559_ (.CLK(net130),
    .D(_00575_),
    .Q(\rbzero.wall_tracer.trackDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20560_ (.CLK(net130),
    .D(_00576_),
    .Q(\rbzero.wall_tracer.trackDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20561_ (.CLK(net136),
    .D(_00577_),
    .Q(\rbzero.wall_tracer.trackDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20562_ (.CLK(net136),
    .D(_00578_),
    .Q(\rbzero.wall_tracer.trackDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20563_ (.CLK(net136),
    .D(_00579_),
    .Q(\rbzero.wall_tracer.trackDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20564_ (.CLK(net123),
    .D(_00580_),
    .Q(\rbzero.wall_tracer.trackDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20565_ (.CLK(net136),
    .D(_00581_),
    .Q(\rbzero.wall_tracer.trackDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20566_ (.CLK(net137),
    .D(_00582_),
    .Q(\rbzero.wall_tracer.trackDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20567_ (.CLK(net137),
    .D(_00583_),
    .Q(\rbzero.wall_tracer.trackDistY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20568_ (.CLK(net137),
    .D(_00584_),
    .Q(\rbzero.wall_tracer.trackDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20569_ (.CLK(net139),
    .D(_00585_),
    .Q(\rbzero.wall_tracer.trackDistY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20570_ (.CLK(net125),
    .D(_00586_),
    .Q(\rbzero.wall_tracer.trackDistY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20571_ (.CLK(net125),
    .D(_00587_),
    .Q(\rbzero.wall_tracer.trackDistY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20572_ (.CLK(net124),
    .D(_00588_),
    .Q(\rbzero.wall_tracer.trackDistY[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20573_ (.CLK(net101),
    .D(_00589_),
    .Q(\rbzero.spi_registers.new_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _20574_ (.CLK(net89),
    .D(_00590_),
    .Q(\rbzero.wall_tracer.rayAddendX[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _20575_ (.CLK(net81),
    .D(_00591_),
    .Q(\rbzero.wall_tracer.rayAddendX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20576_ (.CLK(net81),
    .D(_00592_),
    .Q(\rbzero.wall_tracer.rayAddendX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _20577_ (.CLK(net82),
    .D(_00593_),
    .Q(\rbzero.wall_tracer.rayAddendX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20578_ (.CLK(net89),
    .D(_00594_),
    .Q(\rbzero.wall_tracer.rayAddendX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20579_ (.CLK(net87),
    .D(_00595_),
    .Q(\rbzero.wall_tracer.rayAddendX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20580_ (.CLK(net88),
    .D(_00596_),
    .Q(\rbzero.wall_tracer.rayAddendX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20581_ (.CLK(net93),
    .D(_00597_),
    .Q(\rbzero.wall_tracer.rayAddendX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20582_ (.CLK(net93),
    .D(_00598_),
    .Q(\rbzero.wall_tracer.rayAddendX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20583_ (.CLK(net95),
    .D(_00599_),
    .Q(\rbzero.wall_tracer.rayAddendX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20584_ (.CLK(net95),
    .D(_00600_),
    .Q(\rbzero.wall_tracer.rayAddendX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20585_ (.CLK(net95),
    .D(_00601_),
    .Q(\rbzero.wall_tracer.rayAddendX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20586_ (.CLK(net95),
    .D(_00602_),
    .Q(\rbzero.wall_tracer.rayAddendX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20587_ (.CLK(net90),
    .D(_00603_),
    .Q(\rbzero.wall_tracer.rayAddendX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20588_ (.CLK(net90),
    .D(_00604_),
    .Q(\rbzero.wall_tracer.rayAddendX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20589_ (.CLK(net95),
    .D(_00605_),
    .Q(\rbzero.wall_tracer.rayAddendX[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20590_ (.CLK(net95),
    .D(_00606_),
    .Q(\rbzero.wall_tracer.rayAddendX[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20591_ (.CLK(net96),
    .D(_00607_),
    .Q(\rbzero.map_rom.f4 ));
 sky130_fd_sc_hd__dfxtp_2 _20592_ (.CLK(net97),
    .D(_00608_),
    .Q(\rbzero.map_rom.f3 ));
 sky130_fd_sc_hd__dfxtp_1 _20593_ (.CLK(net97),
    .D(_00609_),
    .Q(\rbzero.map_rom.f2 ));
 sky130_fd_sc_hd__dfxtp_2 _20594_ (.CLK(net92),
    .D(_00610_),
    .Q(\rbzero.map_rom.f1 ));
 sky130_fd_sc_hd__dfxtp_1 _20595_ (.CLK(net96),
    .D(_00611_),
    .Q(\rbzero.map_rom.i_col[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20596_ (.CLK(net80),
    .D(_00612_),
    .Q(\rbzero.wall_tracer.rayAddendY[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _20597_ (.CLK(net80),
    .D(_00613_),
    .Q(\rbzero.wall_tracer.rayAddendY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20598_ (.CLK(net82),
    .D(_00614_),
    .Q(\rbzero.wall_tracer.rayAddendY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _20599_ (.CLK(net82),
    .D(_00615_),
    .Q(\rbzero.wall_tracer.rayAddendY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _20600_ (.CLK(net82),
    .D(_00616_),
    .Q(\rbzero.wall_tracer.rayAddendY[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _20601_ (.CLK(net81),
    .D(_00617_),
    .Q(\rbzero.wall_tracer.rayAddendY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20602_ (.CLK(net82),
    .D(_00618_),
    .Q(\rbzero.wall_tracer.rayAddendY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20603_ (.CLK(net81),
    .D(_00619_),
    .Q(\rbzero.wall_tracer.rayAddendY[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20604_ (.CLK(net81),
    .D(_00620_),
    .Q(\rbzero.wall_tracer.rayAddendY[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20605_ (.CLK(net81),
    .D(_00621_),
    .Q(\rbzero.wall_tracer.rayAddendY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20606_ (.CLK(net90),
    .D(_00622_),
    .Q(\rbzero.wall_tracer.rayAddendY[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20607_ (.CLK(net90),
    .D(_00623_),
    .Q(\rbzero.wall_tracer.rayAddendY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20608_ (.CLK(net90),
    .D(_00624_),
    .Q(\rbzero.wall_tracer.rayAddendY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20609_ (.CLK(net90),
    .D(_00625_),
    .Q(\rbzero.wall_tracer.rayAddendY[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20610_ (.CLK(net92),
    .D(_00626_),
    .Q(\rbzero.wall_tracer.rayAddendY[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20611_ (.CLK(net92),
    .D(_00627_),
    .Q(\rbzero.wall_tracer.rayAddendY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20612_ (.CLK(net92),
    .D(_00628_),
    .Q(\rbzero.wall_tracer.rayAddendY[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20613_ (.CLK(net99),
    .D(_00629_),
    .Q(\rbzero.spi_registers.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20614_ (.CLK(net99),
    .D(_00630_),
    .Q(\rbzero.spi_registers.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20615_ (.CLK(net84),
    .D(_00631_),
    .Q(\rbzero.spi_registers.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20616_ (.CLK(net99),
    .D(_00632_),
    .Q(\rbzero.spi_registers.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20617_ (.CLK(net84),
    .D(_00633_),
    .Q(\rbzero.spi_registers.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20618_ (.CLK(net84),
    .D(_00634_),
    .Q(\rbzero.spi_registers.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20619_ (.CLK(net84),
    .D(_00635_),
    .Q(\rbzero.spi_registers.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20620_ (.CLK(net79),
    .D(_00636_),
    .Q(\rbzero.pov.ready_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20621_ (.CLK(net79),
    .D(_00637_),
    .Q(\rbzero.pov.ready_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20622_ (.CLK(net80),
    .D(_00638_),
    .Q(\rbzero.pov.ready_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20623_ (.CLK(net79),
    .D(_00639_),
    .Q(\rbzero.pov.ready_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20624_ (.CLK(net54),
    .D(_00640_),
    .Q(\rbzero.pov.ready_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20625_ (.CLK(net79),
    .D(_00641_),
    .Q(\rbzero.pov.ready_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20626_ (.CLK(net54),
    .D(_00642_),
    .Q(\rbzero.pov.ready_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20627_ (.CLK(net54),
    .D(_00643_),
    .Q(\rbzero.pov.ready_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20628_ (.CLK(net54),
    .D(_00644_),
    .Q(\rbzero.pov.ready_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20629_ (.CLK(net56),
    .D(_00645_),
    .Q(\rbzero.pov.ready_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20630_ (.CLK(net56),
    .D(_00646_),
    .Q(\rbzero.pov.ready_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20631_ (.CLK(net55),
    .D(_00647_),
    .Q(\rbzero.pov.ready_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20632_ (.CLK(net55),
    .D(_00648_),
    .Q(\rbzero.pov.ready_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20633_ (.CLK(net54),
    .D(_00649_),
    .Q(\rbzero.pov.ready_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20634_ (.CLK(net55),
    .D(_00650_),
    .Q(\rbzero.pov.ready_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20635_ (.CLK(net55),
    .D(_00651_),
    .Q(\rbzero.pov.ready_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20636_ (.CLK(net54),
    .D(_00652_),
    .Q(\rbzero.pov.ready_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20637_ (.CLK(net55),
    .D(_00653_),
    .Q(\rbzero.pov.ready_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20638_ (.CLK(net55),
    .D(_00654_),
    .Q(\rbzero.pov.ready_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20639_ (.CLK(net56),
    .D(_00655_),
    .Q(\rbzero.pov.ready_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20640_ (.CLK(net56),
    .D(_00656_),
    .Q(\rbzero.pov.ready_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20641_ (.CLK(net56),
    .D(_00657_),
    .Q(\rbzero.pov.ready_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20642_ (.CLK(net66),
    .D(_00658_),
    .Q(\rbzero.pov.ready_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20643_ (.CLK(net66),
    .D(_00659_),
    .Q(\rbzero.pov.ready_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20644_ (.CLK(net66),
    .D(_00660_),
    .Q(\rbzero.pov.ready_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20645_ (.CLK(net62),
    .D(_00661_),
    .Q(\rbzero.pov.ready_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20646_ (.CLK(net66),
    .D(_00662_),
    .Q(\rbzero.pov.ready_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20647_ (.CLK(net66),
    .D(_00663_),
    .Q(\rbzero.pov.ready_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20648_ (.CLK(net66),
    .D(_00664_),
    .Q(\rbzero.pov.ready_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20649_ (.CLK(net63),
    .D(_00665_),
    .Q(\rbzero.pov.ready_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20650_ (.CLK(net63),
    .D(_00666_),
    .Q(\rbzero.pov.ready_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20651_ (.CLK(net62),
    .D(_00667_),
    .Q(\rbzero.pov.ready_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20652_ (.CLK(net62),
    .D(_00668_),
    .Q(\rbzero.pov.ready_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _20653_ (.CLK(net62),
    .D(_00669_),
    .Q(\rbzero.pov.ready_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _20654_ (.CLK(net63),
    .D(_00670_),
    .Q(\rbzero.pov.ready_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _20655_ (.CLK(net63),
    .D(_00671_),
    .Q(\rbzero.pov.ready_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _20656_ (.CLK(net63),
    .D(_00672_),
    .Q(\rbzero.pov.ready_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _20657_ (.CLK(net63),
    .D(_00673_),
    .Q(\rbzero.pov.ready_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _20658_ (.CLK(net63),
    .D(_00674_),
    .Q(\rbzero.pov.ready_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _20659_ (.CLK(net60),
    .D(_00675_),
    .Q(\rbzero.pov.ready_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _20660_ (.CLK(net67),
    .D(_00676_),
    .Q(\rbzero.pov.ready_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _20661_ (.CLK(net67),
    .D(_00677_),
    .Q(\rbzero.pov.ready_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _20662_ (.CLK(net67),
    .D(_00678_),
    .Q(\rbzero.pov.ready_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _20663_ (.CLK(net67),
    .D(_00679_),
    .Q(\rbzero.pov.ready_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _20664_ (.CLK(net60),
    .D(_00680_),
    .Q(\rbzero.pov.ready_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _20665_ (.CLK(net60),
    .D(_00681_),
    .Q(\rbzero.pov.ready_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _20666_ (.CLK(net61),
    .D(_00682_),
    .Q(\rbzero.pov.ready_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _20667_ (.CLK(net68),
    .D(_00683_),
    .Q(\rbzero.pov.ready_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _20668_ (.CLK(net78),
    .D(_00684_),
    .Q(\rbzero.pov.ready_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _20669_ (.CLK(net74),
    .D(_00685_),
    .Q(\rbzero.pov.ready_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _20670_ (.CLK(net74),
    .D(_00686_),
    .Q(\rbzero.pov.ready_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _20671_ (.CLK(net74),
    .D(_00687_),
    .Q(\rbzero.pov.ready_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _20672_ (.CLK(net70),
    .D(_00688_),
    .Q(\rbzero.pov.ready_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _20673_ (.CLK(net68),
    .D(_00689_),
    .Q(\rbzero.pov.ready_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _20674_ (.CLK(net68),
    .D(_00690_),
    .Q(\rbzero.pov.ready_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _20675_ (.CLK(net68),
    .D(_00691_),
    .Q(\rbzero.pov.ready_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _20676_ (.CLK(net68),
    .D(_00692_),
    .Q(\rbzero.pov.ready_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _20677_ (.CLK(net67),
    .D(_00693_),
    .Q(\rbzero.pov.ready_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _20678_ (.CLK(net67),
    .D(_00694_),
    .Q(\rbzero.pov.ready_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _20679_ (.CLK(net76),
    .D(_00695_),
    .Q(\rbzero.pov.ready_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _20680_ (.CLK(net74),
    .D(_00696_),
    .Q(\rbzero.pov.ready_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _20681_ (.CLK(net76),
    .D(_00697_),
    .Q(\rbzero.pov.ready_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _20682_ (.CLK(net75),
    .D(_00698_),
    .Q(\rbzero.pov.ready_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _20683_ (.CLK(net76),
    .D(_00699_),
    .Q(\rbzero.pov.ready_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _20684_ (.CLK(net75),
    .D(_00700_),
    .Q(\rbzero.pov.ready_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _20685_ (.CLK(net76),
    .D(_00701_),
    .Q(\rbzero.pov.ready_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _20686_ (.CLK(net76),
    .D(_00702_),
    .Q(\rbzero.pov.ready_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _20687_ (.CLK(net76),
    .D(_00703_),
    .Q(\rbzero.pov.ready_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _20688_ (.CLK(net70),
    .D(_00704_),
    .Q(\rbzero.pov.ready_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _20689_ (.CLK(net71),
    .D(_00705_),
    .Q(\rbzero.pov.ready_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _20690_ (.CLK(net70),
    .D(_00706_),
    .Q(\rbzero.pov.ready_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _20691_ (.CLK(net70),
    .D(_00707_),
    .Q(\rbzero.pov.ready_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _20692_ (.CLK(net70),
    .D(_00708_),
    .Q(\rbzero.pov.ready_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _20693_ (.CLK(net70),
    .D(_00709_),
    .Q(\rbzero.pov.ready_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_2 _20694_ (.CLK(net84),
    .D(_00710_),
    .Q(\rbzero.spi_registers.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20695_ (.CLK(net99),
    .D(_00711_),
    .Q(\rbzero.spi_registers.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20696_ (.CLK(net99),
    .D(_00712_),
    .Q(\rbzero.spi_registers.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20697_ (.CLK(net101),
    .D(_00713_),
    .Q(\rbzero.spi_registers.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20698_ (.CLK(net101),
    .D(_00714_),
    .Q(\rbzero.spi_registers.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20699_ (.CLK(net101),
    .D(_00715_),
    .Q(\rbzero.spi_registers.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20700_ (.CLK(net87),
    .D(_00716_),
    .Q(\rbzero.spi_registers.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20701_ (.CLK(net87),
    .D(_00717_),
    .Q(\rbzero.spi_registers.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20702_ (.CLK(net87),
    .D(_00718_),
    .Q(\rbzero.spi_registers.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20703_ (.CLK(net87),
    .D(_00719_),
    .Q(\rbzero.spi_registers.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20704_ (.CLK(net87),
    .D(_00720_),
    .Q(\rbzero.spi_registers.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20705_ (.CLK(net99),
    .D(_00721_),
    .Q(\rbzero.spi_registers.spi_cmd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20706_ (.CLK(net99),
    .D(_00722_),
    .Q(\rbzero.spi_registers.spi_cmd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20707_ (.CLK(net99),
    .D(_00723_),
    .Q(\rbzero.spi_registers.spi_cmd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20708_ (.CLK(net99),
    .D(_00724_),
    .Q(\rbzero.spi_registers.spi_cmd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20709_ (.CLK(net84),
    .D(_00725_),
    .Q(\rbzero.spi_registers.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20710_ (.CLK(net85),
    .D(_00726_),
    .Q(\rbzero.spi_registers.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _20711_ (.CLK(net109),
    .D(_00727_),
    .Q(\rbzero.spi_registers.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20712_ (.CLK(net99),
    .D(_00728_),
    .Q(\rbzero.spi_registers.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20713_ (.CLK(net109),
    .D(_00729_),
    .Q(\rbzero.spi_registers.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20714_ (.CLK(net85),
    .D(_00730_),
    .Q(\rbzero.spi_registers.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20715_ (.CLK(net85),
    .D(_00731_),
    .Q(\rbzero.spi_registers.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20716_ (.CLK(net93),
    .D(_00732_),
    .Q(\rbzero.otherx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20717_ (.CLK(net93),
    .D(_00733_),
    .Q(\rbzero.otherx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20718_ (.CLK(net93),
    .D(_00734_),
    .Q(\rbzero.otherx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20719_ (.CLK(net88),
    .D(_00735_),
    .Q(\rbzero.otherx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20720_ (.CLK(net93),
    .D(_00736_),
    .Q(\rbzero.otherx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20721_ (.CLK(net93),
    .D(_00737_),
    .Q(\rbzero.othery[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20722_ (.CLK(net101),
    .D(_00738_),
    .Q(\rbzero.othery[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20723_ (.CLK(net93),
    .D(_00739_),
    .Q(\rbzero.othery[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20724_ (.CLK(net94),
    .D(_00740_),
    .Q(\rbzero.othery[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20725_ (.CLK(net101),
    .D(_00741_),
    .Q(\rbzero.othery[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20726_ (.CLK(net101),
    .D(_00742_),
    .Q(\rbzero.row_render.vinf ));
 sky130_fd_sc_hd__dfxtp_1 _20727_ (.CLK(net100),
    .D(_00743_),
    .Q(\rbzero.floor_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20728_ (.CLK(net100),
    .D(_00744_),
    .Q(\rbzero.floor_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20729_ (.CLK(net100),
    .D(_00745_),
    .Q(\rbzero.floor_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20730_ (.CLK(net100),
    .D(_00746_),
    .Q(\rbzero.floor_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20731_ (.CLK(net103),
    .D(_00747_),
    .Q(\rbzero.floor_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20732_ (.CLK(net103),
    .D(_00748_),
    .Q(\rbzero.floor_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20733_ (.CLK(net107),
    .D(_00749_),
    .Q(\rbzero.color_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20734_ (.CLK(net105),
    .D(_00750_),
    .Q(\rbzero.color_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20735_ (.CLK(net107),
    .D(_00751_),
    .Q(\rbzero.color_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20736_ (.CLK(net105),
    .D(_00752_),
    .Q(\rbzero.color_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20737_ (.CLK(net107),
    .D(_00753_),
    .Q(\rbzero.color_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20738_ (.CLK(net105),
    .D(_00754_),
    .Q(\rbzero.color_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20739_ (.CLK(net107),
    .D(_00755_),
    .Q(\rbzero.color_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20740_ (.CLK(net105),
    .D(_00756_),
    .Q(\rbzero.color_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20741_ (.CLK(net107),
    .D(_00757_),
    .Q(\rbzero.color_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20742_ (.CLK(net106),
    .D(_00758_),
    .Q(\rbzero.color_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20743_ (.CLK(net107),
    .D(_00759_),
    .Q(\rbzero.color_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20744_ (.CLK(net105),
    .D(_00760_),
    .Q(\rbzero.color_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20745_ (.CLK(net103),
    .D(_00761_),
    .Q(\rbzero.spi_registers.vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20746_ (.CLK(net103),
    .D(_00762_),
    .Q(\rbzero.spi_registers.vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20747_ (.CLK(net103),
    .D(_00763_),
    .Q(\rbzero.spi_registers.vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20748_ (.CLK(net103),
    .D(_00764_),
    .Q(\rbzero.spi_registers.vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20749_ (.CLK(net104),
    .D(_00765_),
    .Q(\rbzero.spi_registers.vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20750_ (.CLK(net109),
    .D(_00766_),
    .Q(\rbzero.spi_registers.vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20751_ (.CLK(net100),
    .D(_00767_),
    .Q(\rbzero.spi_registers.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _20752_ (.CLK(net105),
    .D(_00768_),
    .Q(\rbzero.spi_registers.new_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20753_ (.CLK(net105),
    .D(_00769_),
    .Q(\rbzero.spi_registers.new_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20754_ (.CLK(net106),
    .D(_00770_),
    .Q(\rbzero.spi_registers.new_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20755_ (.CLK(net106),
    .D(_00771_),
    .Q(\rbzero.spi_registers.new_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20756_ (.CLK(net106),
    .D(_00772_),
    .Q(\rbzero.spi_registers.new_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20757_ (.CLK(net105),
    .D(_00773_),
    .Q(\rbzero.spi_registers.new_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20758_ (.CLK(net106),
    .D(_00774_),
    .Q(\rbzero.spi_registers.got_new_sky ));
 sky130_fd_sc_hd__dfxtp_1 _20759_ (.CLK(net107),
    .D(_00775_),
    .Q(\rbzero.spi_registers.new_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20760_ (.CLK(net105),
    .D(_00776_),
    .Q(\rbzero.spi_registers.new_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20761_ (.CLK(net107),
    .D(_00777_),
    .Q(\rbzero.spi_registers.new_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20762_ (.CLK(net106),
    .D(_00778_),
    .Q(\rbzero.spi_registers.new_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20763_ (.CLK(net107),
    .D(_00779_),
    .Q(\rbzero.spi_registers.new_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20764_ (.CLK(net105),
    .D(_00780_),
    .Q(\rbzero.spi_registers.new_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20765_ (.CLK(net106),
    .D(_00781_),
    .Q(\rbzero.spi_registers.got_new_floor ));
 sky130_fd_sc_hd__dfxtp_1 _20766_ (.CLK(net100),
    .D(_00782_),
    .Q(\rbzero.spi_registers.new_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20767_ (.CLK(net100),
    .D(_00783_),
    .Q(\rbzero.spi_registers.new_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20768_ (.CLK(net100),
    .D(_00784_),
    .Q(\rbzero.spi_registers.new_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20769_ (.CLK(net103),
    .D(_00785_),
    .Q(\rbzero.spi_registers.new_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20770_ (.CLK(net103),
    .D(_00786_),
    .Q(\rbzero.spi_registers.new_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20771_ (.CLK(net103),
    .D(_00787_),
    .Q(\rbzero.spi_registers.new_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20772_ (.CLK(net103),
    .D(_00788_),
    .Q(\rbzero.spi_registers.got_new_leak ));
 sky130_fd_sc_hd__dfxtp_1 _20773_ (.CLK(net87),
    .D(_00789_),
    .Q(\rbzero.spi_registers.new_other[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20774_ (.CLK(net102),
    .D(_00790_),
    .Q(\rbzero.spi_registers.new_other[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20775_ (.CLK(net88),
    .D(_00791_),
    .Q(\rbzero.spi_registers.new_other[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20776_ (.CLK(net88),
    .D(_00792_),
    .Q(\rbzero.spi_registers.new_other[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20777_ (.CLK(net102),
    .D(_00793_),
    .Q(\rbzero.spi_registers.new_other[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20778_ (.CLK(net88),
    .D(_00794_),
    .Q(\rbzero.spi_registers.new_other[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20779_ (.CLK(net88),
    .D(_00795_),
    .Q(\rbzero.spi_registers.new_other[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20780_ (.CLK(net87),
    .D(_00796_),
    .Q(\rbzero.spi_registers.new_other[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20781_ (.CLK(net87),
    .D(_00797_),
    .Q(\rbzero.spi_registers.new_other[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20782_ (.CLK(net88),
    .D(_00798_),
    .Q(\rbzero.spi_registers.new_other[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20783_ (.CLK(net102),
    .D(_00799_),
    .Q(\rbzero.spi_registers.got_new_other ));
 sky130_fd_sc_hd__dfxtp_1 _20784_ (.CLK(net102),
    .D(_00800_),
    .Q(\rbzero.spi_registers.new_vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20785_ (.CLK(net101),
    .D(_00801_),
    .Q(\rbzero.spi_registers.new_vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20786_ (.CLK(net102),
    .D(_00802_),
    .Q(\rbzero.spi_registers.new_vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20787_ (.CLK(net102),
    .D(_00803_),
    .Q(\rbzero.spi_registers.new_vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20788_ (.CLK(net102),
    .D(_00804_),
    .Q(\rbzero.spi_registers.new_vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20789_ (.CLK(net101),
    .D(_00805_),
    .Q(\rbzero.spi_registers.new_vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20790_ (.CLK(net102),
    .D(_00806_),
    .Q(\rbzero.spi_registers.got_new_vshift ));
 sky130_fd_sc_hd__dfxtp_1 _20791_ (.CLK(net91),
    .D(_00807_),
    .Q(\rbzero.pov.ready ));
 sky130_fd_sc_hd__dfxtp_1 _20792_ (.CLK(net84),
    .D(_00808_),
    .Q(\rbzero.pov.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20793_ (.CLK(net86),
    .D(_00809_),
    .Q(\rbzero.pov.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20794_ (.CLK(net84),
    .D(_00810_),
    .Q(\rbzero.pov.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20795_ (.CLK(net84),
    .D(_00811_),
    .Q(\rbzero.pov.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20796_ (.CLK(net84),
    .D(_00812_),
    .Q(\rbzero.pov.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20797_ (.CLK(net86),
    .D(_00813_),
    .Q(\rbzero.pov.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20798_ (.CLK(net86),
    .D(_00814_),
    .Q(\rbzero.pov.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20799_ (.CLK(_00017_),
    .D(_00815_),
    .Q(\rbzero.tex_b0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20800_ (.CLK(_00018_),
    .D(_00816_),
    .Q(\rbzero.tex_b0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20801_ (.CLK(_00019_),
    .D(_00817_),
    .Q(\rbzero.tex_b0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20802_ (.CLK(_00020_),
    .D(_00818_),
    .Q(\rbzero.tex_b0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20803_ (.CLK(_00021_),
    .D(_00819_),
    .Q(\rbzero.tex_b0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20804_ (.CLK(_00022_),
    .D(_00820_),
    .Q(\rbzero.tex_b0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20805_ (.CLK(_00023_),
    .D(_00821_),
    .Q(\rbzero.tex_b0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20806_ (.CLK(_00024_),
    .D(_00822_),
    .Q(\rbzero.tex_b0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20807_ (.CLK(_00025_),
    .D(_00823_),
    .Q(\rbzero.tex_b0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20808_ (.CLK(_00026_),
    .D(_00824_),
    .Q(\rbzero.tex_b0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20809_ (.CLK(_00027_),
    .D(_00825_),
    .Q(\rbzero.tex_b0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20810_ (.CLK(_00028_),
    .D(_00826_),
    .Q(\rbzero.tex_b0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20811_ (.CLK(_00029_),
    .D(_00827_),
    .Q(\rbzero.tex_b0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20812_ (.CLK(_00030_),
    .D(_00828_),
    .Q(\rbzero.tex_b0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20813_ (.CLK(_00031_),
    .D(_00829_),
    .Q(\rbzero.tex_b0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20814_ (.CLK(_00032_),
    .D(_00830_),
    .Q(\rbzero.tex_b0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20815_ (.CLK(_00033_),
    .D(_00831_),
    .Q(\rbzero.tex_b0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20816_ (.CLK(_00034_),
    .D(_00832_),
    .Q(\rbzero.tex_b0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20817_ (.CLK(_00035_),
    .D(_00833_),
    .Q(\rbzero.tex_b0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20818_ (.CLK(_00036_),
    .D(_00834_),
    .Q(\rbzero.tex_b0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20819_ (.CLK(_00037_),
    .D(_00835_),
    .Q(\rbzero.tex_b0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20820_ (.CLK(_00038_),
    .D(_00836_),
    .Q(\rbzero.tex_b0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20821_ (.CLK(_00039_),
    .D(_00837_),
    .Q(\rbzero.tex_b0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20822_ (.CLK(_00040_),
    .D(_00838_),
    .Q(\rbzero.tex_b0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20823_ (.CLK(_00041_),
    .D(_00839_),
    .Q(\rbzero.tex_b0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20824_ (.CLK(_00042_),
    .D(_00840_),
    .Q(\rbzero.tex_b0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20825_ (.CLK(_00043_),
    .D(_00841_),
    .Q(\rbzero.tex_b0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20826_ (.CLK(_00044_),
    .D(_00842_),
    .Q(\rbzero.tex_b0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20827_ (.CLK(_00045_),
    .D(_00843_),
    .Q(\rbzero.tex_b0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20828_ (.CLK(_00046_),
    .D(_00844_),
    .Q(\rbzero.tex_b0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20829_ (.CLK(_00047_),
    .D(_00845_),
    .Q(\rbzero.tex_b0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20830_ (.CLK(_00048_),
    .D(_00846_),
    .Q(\rbzero.tex_b0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20831_ (.CLK(_00049_),
    .D(_00847_),
    .Q(\rbzero.tex_b0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _20832_ (.CLK(_00050_),
    .D(_00848_),
    .Q(\rbzero.tex_b0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _20833_ (.CLK(_00051_),
    .D(_00849_),
    .Q(\rbzero.tex_b0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _20834_ (.CLK(_00052_),
    .D(_00850_),
    .Q(\rbzero.tex_b0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _20835_ (.CLK(_00053_),
    .D(_00851_),
    .Q(\rbzero.tex_b0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _20836_ (.CLK(_00054_),
    .D(_00852_),
    .Q(\rbzero.tex_b0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _20837_ (.CLK(_00055_),
    .D(_00853_),
    .Q(\rbzero.tex_b0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _20838_ (.CLK(_00056_),
    .D(_00854_),
    .Q(\rbzero.tex_b0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _20839_ (.CLK(_00057_),
    .D(_00855_),
    .Q(\rbzero.tex_b0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _20840_ (.CLK(_00058_),
    .D(_00856_),
    .Q(\rbzero.tex_b0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _20841_ (.CLK(_00059_),
    .D(_00857_),
    .Q(\rbzero.tex_b0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _20842_ (.CLK(_00060_),
    .D(_00858_),
    .Q(\rbzero.tex_b0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _20843_ (.CLK(_00061_),
    .D(_00859_),
    .Q(\rbzero.tex_b0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _20844_ (.CLK(_00062_),
    .D(_00860_),
    .Q(\rbzero.tex_b0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _20845_ (.CLK(_00063_),
    .D(_00861_),
    .Q(\rbzero.tex_b0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _20846_ (.CLK(_00064_),
    .D(_00862_),
    .Q(\rbzero.tex_b0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _20847_ (.CLK(_00065_),
    .D(_00863_),
    .Q(\rbzero.tex_b0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _20848_ (.CLK(_00066_),
    .D(_00864_),
    .Q(\rbzero.tex_b0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _20849_ (.CLK(_00067_),
    .D(_00865_),
    .Q(\rbzero.tex_b0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _20850_ (.CLK(_00068_),
    .D(_00866_),
    .Q(\rbzero.tex_b0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _20851_ (.CLK(_00069_),
    .D(_00867_),
    .Q(\rbzero.tex_b0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _20852_ (.CLK(_00070_),
    .D(_00868_),
    .Q(\rbzero.tex_b0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _20853_ (.CLK(_00071_),
    .D(_00869_),
    .Q(\rbzero.tex_b0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _20854_ (.CLK(_00072_),
    .D(_00870_),
    .Q(\rbzero.tex_b0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _20855_ (.CLK(_00073_),
    .D(_00871_),
    .Q(\rbzero.tex_b0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _20856_ (.CLK(_00074_),
    .D(_00872_),
    .Q(\rbzero.tex_b0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _20857_ (.CLK(_00075_),
    .D(_00873_),
    .Q(\rbzero.tex_b0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _20858_ (.CLK(_00076_),
    .D(_00874_),
    .Q(\rbzero.tex_b0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _20859_ (.CLK(_00077_),
    .D(_00875_),
    .Q(\rbzero.tex_b0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _20860_ (.CLK(_00078_),
    .D(_00876_),
    .Q(\rbzero.tex_b0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _20861_ (.CLK(_00079_),
    .D(_00877_),
    .Q(\rbzero.tex_b0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _20862_ (.CLK(_00080_),
    .D(_00878_),
    .Q(\rbzero.tex_b0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _20863_ (.CLK(net79),
    .D(_00879_),
    .Q(\rbzero.pov.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20864_ (.CLK(net79),
    .D(_00880_),
    .Q(\rbzero.pov.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20865_ (.CLK(net79),
    .D(_00881_),
    .Q(\rbzero.pov.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20866_ (.CLK(net79),
    .D(_00882_),
    .Q(\rbzero.pov.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20867_ (.CLK(net79),
    .D(_00883_),
    .Q(\rbzero.pov.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20868_ (.CLK(net54),
    .D(_00884_),
    .Q(\rbzero.pov.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20869_ (.CLK(net54),
    .D(_00885_),
    .Q(\rbzero.pov.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20870_ (.CLK(net54),
    .D(_00886_),
    .Q(\rbzero.pov.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20871_ (.CLK(net54),
    .D(_00887_),
    .Q(\rbzero.pov.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20872_ (.CLK(net59),
    .D(_00888_),
    .Q(\rbzero.pov.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20873_ (.CLK(net56),
    .D(_00889_),
    .Q(\rbzero.pov.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20874_ (.CLK(net58),
    .D(_00890_),
    .Q(\rbzero.pov.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20875_ (.CLK(net58),
    .D(_00891_),
    .Q(\rbzero.pov.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20876_ (.CLK(net58),
    .D(_00892_),
    .Q(\rbzero.pov.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20877_ (.CLK(net55),
    .D(_00893_),
    .Q(\rbzero.pov.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20878_ (.CLK(net58),
    .D(_00894_),
    .Q(\rbzero.pov.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20879_ (.CLK(net59),
    .D(_00895_),
    .Q(\rbzero.pov.spi_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20880_ (.CLK(net58),
    .D(_00896_),
    .Q(\rbzero.pov.spi_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20881_ (.CLK(net55),
    .D(_00897_),
    .Q(\rbzero.pov.spi_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20882_ (.CLK(net58),
    .D(_00898_),
    .Q(\rbzero.pov.spi_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20883_ (.CLK(net58),
    .D(_00899_),
    .Q(\rbzero.pov.spi_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20884_ (.CLK(net58),
    .D(_00900_),
    .Q(\rbzero.pov.spi_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20885_ (.CLK(net56),
    .D(_00901_),
    .Q(\rbzero.pov.spi_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20886_ (.CLK(net66),
    .D(_00902_),
    .Q(\rbzero.pov.spi_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20887_ (.CLK(net62),
    .D(_00903_),
    .Q(\rbzero.pov.spi_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20888_ (.CLK(net62),
    .D(_00904_),
    .Q(\rbzero.pov.spi_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20889_ (.CLK(net64),
    .D(_00905_),
    .Q(\rbzero.pov.spi_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20890_ (.CLK(net66),
    .D(_00906_),
    .Q(\rbzero.pov.spi_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20891_ (.CLK(net64),
    .D(_00907_),
    .Q(\rbzero.pov.spi_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20892_ (.CLK(net62),
    .D(_00908_),
    .Q(\rbzero.pov.spi_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20893_ (.CLK(net62),
    .D(_00909_),
    .Q(\rbzero.pov.spi_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20894_ (.CLK(net62),
    .D(_00910_),
    .Q(\rbzero.pov.spi_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20895_ (.CLK(net62),
    .D(_00911_),
    .Q(\rbzero.pov.spi_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _20896_ (.CLK(net60),
    .D(_00912_),
    .Q(\rbzero.pov.spi_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _20897_ (.CLK(net60),
    .D(_00913_),
    .Q(\rbzero.pov.spi_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _20898_ (.CLK(net60),
    .D(_00914_),
    .Q(\rbzero.pov.spi_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _20899_ (.CLK(net60),
    .D(_00915_),
    .Q(\rbzero.pov.spi_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _20900_ (.CLK(net60),
    .D(_00916_),
    .Q(\rbzero.pov.spi_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _20901_ (.CLK(net60),
    .D(_00917_),
    .Q(\rbzero.pov.spi_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _20902_ (.CLK(net60),
    .D(_00918_),
    .Q(\rbzero.pov.spi_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _20903_ (.CLK(net61),
    .D(_00919_),
    .Q(\rbzero.pov.spi_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _20904_ (.CLK(net67),
    .D(_00920_),
    .Q(\rbzero.pov.spi_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _20905_ (.CLK(net67),
    .D(_00921_),
    .Q(\rbzero.pov.spi_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _20906_ (.CLK(net61),
    .D(_00922_),
    .Q(\rbzero.pov.spi_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _20907_ (.CLK(net61),
    .D(_00923_),
    .Q(\rbzero.pov.spi_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _20908_ (.CLK(net61),
    .D(_00924_),
    .Q(\rbzero.pov.spi_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _20909_ (.CLK(net61),
    .D(_00925_),
    .Q(\rbzero.pov.spi_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _20910_ (.CLK(net61),
    .D(_00926_),
    .Q(\rbzero.pov.spi_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _20911_ (.CLK(net78),
    .D(_00927_),
    .Q(\rbzero.pov.spi_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _20912_ (.CLK(net78),
    .D(_00928_),
    .Q(\rbzero.pov.spi_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _20913_ (.CLK(net78),
    .D(_00929_),
    .Q(\rbzero.pov.spi_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _20914_ (.CLK(net74),
    .D(_00930_),
    .Q(\rbzero.pov.spi_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _20915_ (.CLK(net68),
    .D(_00931_),
    .Q(\rbzero.pov.spi_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _20916_ (.CLK(net69),
    .D(_00932_),
    .Q(\rbzero.pov.spi_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _20917_ (.CLK(net68),
    .D(_00933_),
    .Q(\rbzero.pov.spi_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _20918_ (.CLK(net68),
    .D(_00934_),
    .Q(\rbzero.pov.spi_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _20919_ (.CLK(net68),
    .D(_00935_),
    .Q(\rbzero.pov.spi_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _20920_ (.CLK(net67),
    .D(_00936_),
    .Q(\rbzero.pov.spi_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _20921_ (.CLK(net68),
    .D(_00937_),
    .Q(\rbzero.pov.spi_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _20922_ (.CLK(net74),
    .D(_00938_),
    .Q(\rbzero.pov.spi_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _20923_ (.CLK(net74),
    .D(_00939_),
    .Q(\rbzero.pov.spi_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _20924_ (.CLK(net75),
    .D(_00940_),
    .Q(\rbzero.pov.spi_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _20925_ (.CLK(net75),
    .D(_00941_),
    .Q(\rbzero.pov.spi_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _20926_ (.CLK(net75),
    .D(_00942_),
    .Q(\rbzero.pov.spi_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _20927_ (.CLK(net75),
    .D(_00943_),
    .Q(\rbzero.pov.spi_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _20928_ (.CLK(net75),
    .D(_00944_),
    .Q(\rbzero.pov.spi_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _20929_ (.CLK(net74),
    .D(_00945_),
    .Q(\rbzero.pov.spi_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _20930_ (.CLK(net74),
    .D(_00946_),
    .Q(\rbzero.pov.spi_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _20931_ (.CLK(net74),
    .D(_00947_),
    .Q(\rbzero.pov.spi_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _20932_ (.CLK(net67),
    .D(_00948_),
    .Q(\rbzero.pov.spi_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _20933_ (.CLK(net69),
    .D(_00949_),
    .Q(\rbzero.pov.spi_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _20934_ (.CLK(net69),
    .D(_00950_),
    .Q(\rbzero.pov.spi_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _20935_ (.CLK(net69),
    .D(_00951_),
    .Q(\rbzero.pov.spi_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _20936_ (.CLK(net70),
    .D(_00952_),
    .Q(\rbzero.pov.spi_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _20937_ (.CLK(net93),
    .D(_00953_),
    .Q(\rbzero.pov.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20938_ (.CLK(net87),
    .D(_00954_),
    .Q(\rbzero.pov.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _20939_ (.CLK(net100),
    .D(_00955_),
    .Q(\rbzero.pov.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20940_ (.CLK(net85),
    .D(_00956_),
    .Q(\rbzero.pov.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20941_ (.CLK(net104),
    .D(_00957_),
    .Q(\rbzero.pov.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20942_ (.CLK(net85),
    .D(_00958_),
    .Q(\rbzero.pov.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20943_ (.CLK(net85),
    .D(_00959_),
    .Q(\rbzero.pov.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_4 _20944_ (.CLK(net76),
    .D(_00960_),
    .Q(\rbzero.debug_overlay.playerX[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _20945_ (.CLK(net77),
    .D(_00961_),
    .Q(\rbzero.debug_overlay.playerX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20946_ (.CLK(net77),
    .D(_00962_),
    .Q(\rbzero.debug_overlay.playerX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20947_ (.CLK(net116),
    .D(_00963_),
    .Q(\rbzero.debug_overlay.playerX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20948_ (.CLK(net77),
    .D(_00964_),
    .Q(\rbzero.debug_overlay.playerX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20949_ (.CLK(net116),
    .D(_00965_),
    .Q(\rbzero.debug_overlay.playerX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20950_ (.CLK(net76),
    .D(_00966_),
    .Q(\rbzero.debug_overlay.playerX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _20951_ (.CLK(net76),
    .D(_00967_),
    .Q(\rbzero.debug_overlay.playerX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20952_ (.CLK(net116),
    .D(_00968_),
    .Q(\rbzero.debug_overlay.playerX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20953_ (.CLK(net91),
    .D(_00969_),
    .Q(\rbzero.debug_overlay.playerX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20954_ (.CLK(net71),
    .D(_00970_),
    .Q(\rbzero.debug_overlay.playerX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20955_ (.CLK(net91),
    .D(_00971_),
    .Q(\rbzero.debug_overlay.playerX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20956_ (.CLK(net91),
    .D(_00972_),
    .Q(\rbzero.debug_overlay.playerX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20957_ (.CLK(net70),
    .D(_00973_),
    .Q(\rbzero.debug_overlay.playerX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20958_ (.CLK(net70),
    .D(_00974_),
    .Q(\rbzero.debug_overlay.playerX[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20959_ (.CLK(net91),
    .D(_00975_),
    .Q(\rbzero.debug_overlay.playerY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _20960_ (.CLK(net91),
    .D(_00976_),
    .Q(\rbzero.debug_overlay.playerY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20961_ (.CLK(net91),
    .D(_00977_),
    .Q(\rbzero.debug_overlay.playerY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20962_ (.CLK(net91),
    .D(_00978_),
    .Q(\rbzero.debug_overlay.playerY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20963_ (.CLK(net116),
    .D(_00979_),
    .Q(\rbzero.debug_overlay.playerY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20964_ (.CLK(net116),
    .D(_00980_),
    .Q(\rbzero.debug_overlay.playerY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20965_ (.CLK(net76),
    .D(_00981_),
    .Q(\rbzero.debug_overlay.playerY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _20966_ (.CLK(net116),
    .D(_00982_),
    .Q(\rbzero.debug_overlay.playerY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20967_ (.CLK(net91),
    .D(_00983_),
    .Q(\rbzero.debug_overlay.playerY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20968_ (.CLK(net71),
    .D(_00984_),
    .Q(\rbzero.debug_overlay.playerY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20969_ (.CLK(net71),
    .D(_00985_),
    .Q(\rbzero.debug_overlay.playerY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20970_ (.CLK(net71),
    .D(_00986_),
    .Q(\rbzero.debug_overlay.playerY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20971_ (.CLK(net71),
    .D(_00987_),
    .Q(\rbzero.debug_overlay.playerY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20972_ (.CLK(net70),
    .D(_00988_),
    .Q(\rbzero.debug_overlay.playerY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20973_ (.CLK(net91),
    .D(_00989_),
    .Q(\rbzero.debug_overlay.playerY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20974_ (.CLK(net63),
    .D(_00990_),
    .Q(\rbzero.debug_overlay.facingX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20975_ (.CLK(net90),
    .D(_00991_),
    .Q(\rbzero.debug_overlay.facingX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20976_ (.CLK(net63),
    .D(_00992_),
    .Q(\rbzero.debug_overlay.facingX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20977_ (.CLK(net63),
    .D(_00993_),
    .Q(\rbzero.debug_overlay.facingX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20978_ (.CLK(net64),
    .D(_00994_),
    .Q(\rbzero.debug_overlay.facingX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20979_ (.CLK(net65),
    .D(_00995_),
    .Q(\rbzero.debug_overlay.facingX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20980_ (.CLK(net90),
    .D(_00996_),
    .Q(\rbzero.debug_overlay.facingX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20981_ (.CLK(net90),
    .D(_00997_),
    .Q(\rbzero.debug_overlay.facingX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20982_ (.CLK(net65),
    .D(_00998_),
    .Q(\rbzero.debug_overlay.facingX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20983_ (.CLK(net65),
    .D(_00999_),
    .Q(\rbzero.debug_overlay.facingX[0] ));
 sky130_fd_sc_hd__dfxtp_4 _20984_ (.CLK(net65),
    .D(_01000_),
    .Q(\rbzero.debug_overlay.facingX[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20985_ (.CLK(net65),
    .D(_01001_),
    .Q(\rbzero.debug_overlay.facingY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20986_ (.CLK(net65),
    .D(_01002_),
    .Q(\rbzero.debug_overlay.facingY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20987_ (.CLK(net65),
    .D(_01003_),
    .Q(\rbzero.debug_overlay.facingY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20988_ (.CLK(net65),
    .D(_01004_),
    .Q(\rbzero.debug_overlay.facingY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20989_ (.CLK(net65),
    .D(_01005_),
    .Q(\rbzero.debug_overlay.facingY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20990_ (.CLK(net66),
    .D(_01006_),
    .Q(\rbzero.debug_overlay.facingY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20991_ (.CLK(net90),
    .D(_01007_),
    .Q(\rbzero.debug_overlay.facingY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _20992_ (.CLK(net65),
    .D(_01008_),
    .Q(\rbzero.debug_overlay.facingY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20993_ (.CLK(net72),
    .D(_01009_),
    .Q(\rbzero.debug_overlay.facingY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20994_ (.CLK(net56),
    .D(_01010_),
    .Q(\rbzero.debug_overlay.facingY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20995_ (.CLK(net66),
    .D(_01011_),
    .Q(\rbzero.debug_overlay.facingY[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20996_ (.CLK(net55),
    .D(_01012_),
    .Q(\rbzero.debug_overlay.vplaneX[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _20997_ (.CLK(net56),
    .D(_01013_),
    .Q(\rbzero.debug_overlay.vplaneX[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _20998_ (.CLK(net59),
    .D(_01014_),
    .Q(\rbzero.debug_overlay.vplaneX[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _20999_ (.CLK(net55),
    .D(_01015_),
    .Q(\rbzero.debug_overlay.vplaneX[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21000_ (.CLK(net57),
    .D(_01016_),
    .Q(\rbzero.debug_overlay.vplaneX[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _21001_ (.CLK(net81),
    .D(_01017_),
    .Q(\rbzero.debug_overlay.vplaneX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21002_ (.CLK(net57),
    .D(_01018_),
    .Q(\rbzero.debug_overlay.vplaneX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21003_ (.CLK(net57),
    .D(_01019_),
    .Q(\rbzero.debug_overlay.vplaneX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21004_ (.CLK(net82),
    .D(_01020_),
    .Q(\rbzero.debug_overlay.vplaneX[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21005_ (.CLK(net56),
    .D(_01021_),
    .Q(\rbzero.debug_overlay.vplaneX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21006_ (.CLK(net82),
    .D(_01022_),
    .Q(\rbzero.debug_overlay.vplaneX[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21007_ (.CLK(net79),
    .D(_01023_),
    .Q(\rbzero.debug_overlay.vplaneY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21008_ (.CLK(net80),
    .D(_01024_),
    .Q(\rbzero.debug_overlay.vplaneY[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _21009_ (.CLK(net80),
    .D(_01025_),
    .Q(\rbzero.debug_overlay.vplaneY[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _21010_ (.CLK(net80),
    .D(_01026_),
    .Q(\rbzero.debug_overlay.vplaneY[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21011_ (.CLK(net81),
    .D(_01027_),
    .Q(\rbzero.debug_overlay.vplaneY[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _21012_ (.CLK(net80),
    .D(_01028_),
    .Q(\rbzero.debug_overlay.vplaneY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21013_ (.CLK(net80),
    .D(_01029_),
    .Q(\rbzero.debug_overlay.vplaneY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21014_ (.CLK(net81),
    .D(_01030_),
    .Q(\rbzero.debug_overlay.vplaneY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21015_ (.CLK(net57),
    .D(_01031_),
    .Q(\rbzero.debug_overlay.vplaneY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21016_ (.CLK(net57),
    .D(_01032_),
    .Q(\rbzero.debug_overlay.vplaneY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21017_ (.CLK(net81),
    .D(_01033_),
    .Q(\rbzero.debug_overlay.vplaneY[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21018_ (.CLK(net80),
    .D(_01034_),
    .Q(\rbzero.pov.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _21019_ (.CLK(net94),
    .D(_01035_),
    .Q(\rbzero.vga_sync.vsync ));
 sky130_fd_sc_hd__dfxtp_1 _21020_ (.CLK(net94),
    .D(_01036_),
    .Q(\rbzero.hsync ));
 sky130_fd_sc_hd__dfxtp_1 _21021_ (.CLK(net110),
    .D(_01037_),
    .Q(\gpout0.vpos[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21022_ (.CLK(net110),
    .D(_01038_),
    .Q(\gpout0.vpos[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21023_ (.CLK(net110),
    .D(_01039_),
    .Q(\gpout0.vpos[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21024_ (.CLK(net109),
    .D(_01040_),
    .Q(\gpout0.vpos[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21025_ (.CLK(net95),
    .D(_01041_),
    .Q(\gpout0.vpos[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21026_ (.CLK(net93),
    .D(_01042_),
    .Q(\gpout0.vpos[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21027_ (.CLK(net109),
    .D(_01043_),
    .Q(\gpout0.vpos[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21028_ (.CLK(net110),
    .D(_01044_),
    .Q(\gpout0.vpos[7] ));
 sky130_fd_sc_hd__dfxtp_2 _21029_ (.CLK(net109),
    .D(_01045_),
    .Q(\gpout0.vpos[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21030_ (.CLK(net110),
    .D(_01046_),
    .Q(\gpout0.vpos[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21031_ (.CLK(net101),
    .D(_01047_),
    .Q(\rbzero.spi_registers.got_new_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21032_ (.CLK(_00081_),
    .D(_01048_),
    .Q(\rbzero.tex_g0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21033_ (.CLK(_00082_),
    .D(_01049_),
    .Q(\rbzero.tex_g0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21034_ (.CLK(_00083_),
    .D(_01050_),
    .Q(\rbzero.tex_g0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21035_ (.CLK(_00084_),
    .D(_01051_),
    .Q(\rbzero.tex_g0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21036_ (.CLK(_00085_),
    .D(_01052_),
    .Q(\rbzero.tex_g0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21037_ (.CLK(_00086_),
    .D(_01053_),
    .Q(\rbzero.tex_g0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21038_ (.CLK(_00087_),
    .D(_01054_),
    .Q(\rbzero.tex_g0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21039_ (.CLK(_00088_),
    .D(_01055_),
    .Q(\rbzero.tex_g0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21040_ (.CLK(_00089_),
    .D(_01056_),
    .Q(\rbzero.tex_g0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21041_ (.CLK(_00090_),
    .D(_01057_),
    .Q(\rbzero.tex_g0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21042_ (.CLK(_00091_),
    .D(_01058_),
    .Q(\rbzero.tex_g0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21043_ (.CLK(_00092_),
    .D(_01059_),
    .Q(\rbzero.tex_g0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21044_ (.CLK(_00093_),
    .D(_01060_),
    .Q(\rbzero.tex_g0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21045_ (.CLK(_00094_),
    .D(_01061_),
    .Q(\rbzero.tex_g0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21046_ (.CLK(_00095_),
    .D(_01062_),
    .Q(\rbzero.tex_g0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21047_ (.CLK(_00096_),
    .D(_01063_),
    .Q(\rbzero.tex_g0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21048_ (.CLK(_00097_),
    .D(_01064_),
    .Q(\rbzero.tex_g0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21049_ (.CLK(_00098_),
    .D(_01065_),
    .Q(\rbzero.tex_g0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21050_ (.CLK(_00099_),
    .D(_01066_),
    .Q(\rbzero.tex_g0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21051_ (.CLK(_00100_),
    .D(_01067_),
    .Q(\rbzero.tex_g0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21052_ (.CLK(_00101_),
    .D(_01068_),
    .Q(\rbzero.tex_g0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21053_ (.CLK(_00102_),
    .D(_01069_),
    .Q(\rbzero.tex_g0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21054_ (.CLK(_00103_),
    .D(_01070_),
    .Q(\rbzero.tex_g0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21055_ (.CLK(_00104_),
    .D(_01071_),
    .Q(\rbzero.tex_g0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21056_ (.CLK(_00105_),
    .D(_01072_),
    .Q(\rbzero.tex_g0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21057_ (.CLK(_00106_),
    .D(_01073_),
    .Q(\rbzero.tex_g0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21058_ (.CLK(_00107_),
    .D(_01074_),
    .Q(\rbzero.tex_g0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21059_ (.CLK(_00108_),
    .D(_01075_),
    .Q(\rbzero.tex_g0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21060_ (.CLK(_00109_),
    .D(_01076_),
    .Q(\rbzero.tex_g0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21061_ (.CLK(_00110_),
    .D(_01077_),
    .Q(\rbzero.tex_g0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21062_ (.CLK(_00111_),
    .D(_01078_),
    .Q(\rbzero.tex_g0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21063_ (.CLK(_00112_),
    .D(_01079_),
    .Q(\rbzero.tex_g0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21064_ (.CLK(_00113_),
    .D(_01080_),
    .Q(\rbzero.tex_g0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21065_ (.CLK(_00114_),
    .D(_01081_),
    .Q(\rbzero.tex_g0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21066_ (.CLK(_00115_),
    .D(_01082_),
    .Q(\rbzero.tex_g0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21067_ (.CLK(_00116_),
    .D(_01083_),
    .Q(\rbzero.tex_g0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21068_ (.CLK(_00117_),
    .D(_01084_),
    .Q(\rbzero.tex_g0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21069_ (.CLK(_00118_),
    .D(_01085_),
    .Q(\rbzero.tex_g0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21070_ (.CLK(_00119_),
    .D(_01086_),
    .Q(\rbzero.tex_g0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21071_ (.CLK(_00120_),
    .D(_01087_),
    .Q(\rbzero.tex_g0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21072_ (.CLK(_00121_),
    .D(_01088_),
    .Q(\rbzero.tex_g0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21073_ (.CLK(_00122_),
    .D(_01089_),
    .Q(\rbzero.tex_g0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21074_ (.CLK(_00123_),
    .D(_01090_),
    .Q(\rbzero.tex_g0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21075_ (.CLK(_00124_),
    .D(_01091_),
    .Q(\rbzero.tex_g0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21076_ (.CLK(_00125_),
    .D(_01092_),
    .Q(\rbzero.tex_g0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21077_ (.CLK(_00126_),
    .D(_01093_),
    .Q(\rbzero.tex_g0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21078_ (.CLK(_00127_),
    .D(_01094_),
    .Q(\rbzero.tex_g0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21079_ (.CLK(_00128_),
    .D(_01095_),
    .Q(\rbzero.tex_g0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21080_ (.CLK(_00129_),
    .D(_01096_),
    .Q(\rbzero.tex_g0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21081_ (.CLK(_00130_),
    .D(_01097_),
    .Q(\rbzero.tex_g0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21082_ (.CLK(_00131_),
    .D(_01098_),
    .Q(\rbzero.tex_g0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21083_ (.CLK(_00132_),
    .D(_01099_),
    .Q(\rbzero.tex_g0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21084_ (.CLK(_00133_),
    .D(_01100_),
    .Q(\rbzero.tex_g0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21085_ (.CLK(_00134_),
    .D(_01101_),
    .Q(\rbzero.tex_g0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21086_ (.CLK(_00135_),
    .D(_01102_),
    .Q(\rbzero.tex_g0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21087_ (.CLK(_00136_),
    .D(_01103_),
    .Q(\rbzero.tex_g0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21088_ (.CLK(_00137_),
    .D(_01104_),
    .Q(\rbzero.tex_g0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21089_ (.CLK(_00138_),
    .D(_01105_),
    .Q(\rbzero.tex_g0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21090_ (.CLK(_00139_),
    .D(_01106_),
    .Q(\rbzero.tex_g0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21091_ (.CLK(_00140_),
    .D(_01107_),
    .Q(\rbzero.tex_g0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21092_ (.CLK(_00141_),
    .D(_01108_),
    .Q(\rbzero.tex_g0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21093_ (.CLK(_00142_),
    .D(_01109_),
    .Q(\rbzero.tex_g0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21094_ (.CLK(_00143_),
    .D(_01110_),
    .Q(\rbzero.tex_g0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21095_ (.CLK(_00144_),
    .D(_01111_),
    .Q(\rbzero.tex_g0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21096_ (.CLK(_00145_),
    .D(_01112_),
    .Q(\rbzero.tex_g1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21097_ (.CLK(_00146_),
    .D(_01113_),
    .Q(\rbzero.tex_g1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21098_ (.CLK(_00147_),
    .D(_01114_),
    .Q(\rbzero.tex_g1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21099_ (.CLK(_00148_),
    .D(_01115_),
    .Q(\rbzero.tex_g1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21100_ (.CLK(_00149_),
    .D(_01116_),
    .Q(\rbzero.tex_g1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21101_ (.CLK(_00150_),
    .D(_01117_),
    .Q(\rbzero.tex_g1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21102_ (.CLK(_00151_),
    .D(_01118_),
    .Q(\rbzero.tex_g1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21103_ (.CLK(_00152_),
    .D(_01119_),
    .Q(\rbzero.tex_g1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21104_ (.CLK(_00153_),
    .D(_01120_),
    .Q(\rbzero.tex_g1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21105_ (.CLK(_00154_),
    .D(_01121_),
    .Q(\rbzero.tex_g1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21106_ (.CLK(_00155_),
    .D(_01122_),
    .Q(\rbzero.tex_g1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21107_ (.CLK(_00156_),
    .D(_01123_),
    .Q(\rbzero.tex_g1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21108_ (.CLK(_00157_),
    .D(_01124_),
    .Q(\rbzero.tex_g1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21109_ (.CLK(_00158_),
    .D(_01125_),
    .Q(\rbzero.tex_g1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21110_ (.CLK(_00159_),
    .D(_01126_),
    .Q(\rbzero.tex_g1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21111_ (.CLK(_00160_),
    .D(_01127_),
    .Q(\rbzero.tex_g1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21112_ (.CLK(_00161_),
    .D(_01128_),
    .Q(\rbzero.tex_g1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21113_ (.CLK(_00162_),
    .D(_01129_),
    .Q(\rbzero.tex_g1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21114_ (.CLK(_00163_),
    .D(_01130_),
    .Q(\rbzero.tex_g1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21115_ (.CLK(_00164_),
    .D(_01131_),
    .Q(\rbzero.tex_g1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21116_ (.CLK(_00165_),
    .D(_01132_),
    .Q(\rbzero.tex_g1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21117_ (.CLK(_00166_),
    .D(_01133_),
    .Q(\rbzero.tex_g1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21118_ (.CLK(_00167_),
    .D(_01134_),
    .Q(\rbzero.tex_g1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21119_ (.CLK(_00168_),
    .D(_01135_),
    .Q(\rbzero.tex_g1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21120_ (.CLK(_00169_),
    .D(_01136_),
    .Q(\rbzero.tex_g1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21121_ (.CLK(_00170_),
    .D(_01137_),
    .Q(\rbzero.tex_g1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21122_ (.CLK(_00171_),
    .D(_01138_),
    .Q(\rbzero.tex_g1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21123_ (.CLK(_00172_),
    .D(_01139_),
    .Q(\rbzero.tex_g1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21124_ (.CLK(_00173_),
    .D(_01140_),
    .Q(\rbzero.tex_g1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21125_ (.CLK(_00174_),
    .D(_01141_),
    .Q(\rbzero.tex_g1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21126_ (.CLK(_00175_),
    .D(_01142_),
    .Q(\rbzero.tex_g1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21127_ (.CLK(_00176_),
    .D(_01143_),
    .Q(\rbzero.tex_g1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21128_ (.CLK(_00177_),
    .D(_01144_),
    .Q(\rbzero.tex_g1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21129_ (.CLK(_00178_),
    .D(_01145_),
    .Q(\rbzero.tex_g1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21130_ (.CLK(_00179_),
    .D(_01146_),
    .Q(\rbzero.tex_g1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21131_ (.CLK(_00180_),
    .D(_01147_),
    .Q(\rbzero.tex_g1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21132_ (.CLK(_00181_),
    .D(_01148_),
    .Q(\rbzero.tex_g1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21133_ (.CLK(_00182_),
    .D(_01149_),
    .Q(\rbzero.tex_g1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21134_ (.CLK(_00183_),
    .D(_01150_),
    .Q(\rbzero.tex_g1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21135_ (.CLK(_00184_),
    .D(_01151_),
    .Q(\rbzero.tex_g1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21136_ (.CLK(_00185_),
    .D(_01152_),
    .Q(\rbzero.tex_g1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21137_ (.CLK(_00186_),
    .D(_01153_),
    .Q(\rbzero.tex_g1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21138_ (.CLK(_00187_),
    .D(_01154_),
    .Q(\rbzero.tex_g1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21139_ (.CLK(_00188_),
    .D(_01155_),
    .Q(\rbzero.tex_g1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21140_ (.CLK(_00189_),
    .D(_01156_),
    .Q(\rbzero.tex_g1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21141_ (.CLK(_00190_),
    .D(_01157_),
    .Q(\rbzero.tex_g1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21142_ (.CLK(_00191_),
    .D(_01158_),
    .Q(\rbzero.tex_g1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21143_ (.CLK(_00192_),
    .D(_01159_),
    .Q(\rbzero.tex_g1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21144_ (.CLK(_00193_),
    .D(_01160_),
    .Q(\rbzero.tex_g1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21145_ (.CLK(_00194_),
    .D(_01161_),
    .Q(\rbzero.tex_g1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21146_ (.CLK(_00195_),
    .D(_01162_),
    .Q(\rbzero.tex_g1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21147_ (.CLK(_00196_),
    .D(_01163_),
    .Q(\rbzero.tex_g1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21148_ (.CLK(_00197_),
    .D(_01164_),
    .Q(\rbzero.tex_g1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21149_ (.CLK(_00198_),
    .D(_01165_),
    .Q(\rbzero.tex_g1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21150_ (.CLK(_00199_),
    .D(_01166_),
    .Q(\rbzero.tex_g1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21151_ (.CLK(_00200_),
    .D(_01167_),
    .Q(\rbzero.tex_g1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21152_ (.CLK(_00201_),
    .D(_01168_),
    .Q(\rbzero.tex_g1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21153_ (.CLK(_00202_),
    .D(_01169_),
    .Q(\rbzero.tex_g1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21154_ (.CLK(_00203_),
    .D(_01170_),
    .Q(\rbzero.tex_g1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21155_ (.CLK(_00204_),
    .D(_01171_),
    .Q(\rbzero.tex_g1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21156_ (.CLK(_00205_),
    .D(_01172_),
    .Q(\rbzero.tex_g1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21157_ (.CLK(_00206_),
    .D(_01173_),
    .Q(\rbzero.tex_g1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21158_ (.CLK(_00207_),
    .D(_01174_),
    .Q(\rbzero.tex_g1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21159_ (.CLK(_00208_),
    .D(_01175_),
    .Q(\rbzero.tex_g1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21160_ (.CLK(_00209_),
    .D(_01176_),
    .Q(\rbzero.tex_r0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21161_ (.CLK(_00210_),
    .D(_01177_),
    .Q(\rbzero.tex_r0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21162_ (.CLK(_00211_),
    .D(_01178_),
    .Q(\rbzero.tex_r0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21163_ (.CLK(_00212_),
    .D(_01179_),
    .Q(\rbzero.tex_r0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21164_ (.CLK(_00213_),
    .D(_01180_),
    .Q(\rbzero.tex_r0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21165_ (.CLK(_00214_),
    .D(_01181_),
    .Q(\rbzero.tex_r0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21166_ (.CLK(_00215_),
    .D(_01182_),
    .Q(\rbzero.tex_r0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21167_ (.CLK(_00216_),
    .D(_01183_),
    .Q(\rbzero.tex_r0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21168_ (.CLK(_00217_),
    .D(_01184_),
    .Q(\rbzero.tex_r0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21169_ (.CLK(_00218_),
    .D(_01185_),
    .Q(\rbzero.tex_r0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21170_ (.CLK(_00219_),
    .D(_01186_),
    .Q(\rbzero.tex_r0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21171_ (.CLK(_00220_),
    .D(_01187_),
    .Q(\rbzero.tex_r0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21172_ (.CLK(_00221_),
    .D(_01188_),
    .Q(\rbzero.tex_r0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21173_ (.CLK(_00222_),
    .D(_01189_),
    .Q(\rbzero.tex_r0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21174_ (.CLK(_00223_),
    .D(_01190_),
    .Q(\rbzero.tex_r0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21175_ (.CLK(_00224_),
    .D(_01191_),
    .Q(\rbzero.tex_r0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21176_ (.CLK(_00225_),
    .D(_01192_),
    .Q(\rbzero.tex_r0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21177_ (.CLK(_00226_),
    .D(_01193_),
    .Q(\rbzero.tex_r0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21178_ (.CLK(_00227_),
    .D(_01194_),
    .Q(\rbzero.tex_r0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21179_ (.CLK(_00228_),
    .D(_01195_),
    .Q(\rbzero.tex_r0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21180_ (.CLK(_00229_),
    .D(_01196_),
    .Q(\rbzero.tex_r0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21181_ (.CLK(_00230_),
    .D(_01197_),
    .Q(\rbzero.tex_r0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21182_ (.CLK(_00231_),
    .D(_01198_),
    .Q(\rbzero.tex_r0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21183_ (.CLK(_00232_),
    .D(_01199_),
    .Q(\rbzero.tex_r0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21184_ (.CLK(_00233_),
    .D(_01200_),
    .Q(\rbzero.tex_r0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21185_ (.CLK(_00234_),
    .D(_01201_),
    .Q(\rbzero.tex_r0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21186_ (.CLK(_00235_),
    .D(_01202_),
    .Q(\rbzero.tex_r0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21187_ (.CLK(_00236_),
    .D(_01203_),
    .Q(\rbzero.tex_r0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21188_ (.CLK(_00237_),
    .D(_01204_),
    .Q(\rbzero.tex_r0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21189_ (.CLK(_00238_),
    .D(_01205_),
    .Q(\rbzero.tex_r0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21190_ (.CLK(_00239_),
    .D(_01206_),
    .Q(\rbzero.tex_r0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21191_ (.CLK(_00240_),
    .D(_01207_),
    .Q(\rbzero.tex_r0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21192_ (.CLK(_00241_),
    .D(_01208_),
    .Q(\rbzero.tex_r0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21193_ (.CLK(_00242_),
    .D(_01209_),
    .Q(\rbzero.tex_r0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21194_ (.CLK(_00243_),
    .D(_01210_),
    .Q(\rbzero.tex_r0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21195_ (.CLK(_00244_),
    .D(_01211_),
    .Q(\rbzero.tex_r0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21196_ (.CLK(_00245_),
    .D(_01212_),
    .Q(\rbzero.tex_r0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21197_ (.CLK(_00246_),
    .D(_01213_),
    .Q(\rbzero.tex_r0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21198_ (.CLK(_00247_),
    .D(_01214_),
    .Q(\rbzero.tex_r0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21199_ (.CLK(_00248_),
    .D(_01215_),
    .Q(\rbzero.tex_r0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21200_ (.CLK(_00249_),
    .D(_01216_),
    .Q(\rbzero.tex_r0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21201_ (.CLK(_00250_),
    .D(_01217_),
    .Q(\rbzero.tex_r0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21202_ (.CLK(_00251_),
    .D(_01218_),
    .Q(\rbzero.tex_r0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21203_ (.CLK(_00252_),
    .D(_01219_),
    .Q(\rbzero.tex_r0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21204_ (.CLK(_00253_),
    .D(_01220_),
    .Q(\rbzero.tex_r0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21205_ (.CLK(_00254_),
    .D(_01221_),
    .Q(\rbzero.tex_r0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21206_ (.CLK(_00255_),
    .D(_01222_),
    .Q(\rbzero.tex_r0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21207_ (.CLK(_00256_),
    .D(_01223_),
    .Q(\rbzero.tex_r0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21208_ (.CLK(_00257_),
    .D(_01224_),
    .Q(\rbzero.tex_r0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21209_ (.CLK(_00258_),
    .D(_01225_),
    .Q(\rbzero.tex_r0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21210_ (.CLK(_00259_),
    .D(_01226_),
    .Q(\rbzero.tex_r0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21211_ (.CLK(_00260_),
    .D(_01227_),
    .Q(\rbzero.tex_r0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21212_ (.CLK(_00261_),
    .D(_01228_),
    .Q(\rbzero.tex_r0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21213_ (.CLK(_00262_),
    .D(_01229_),
    .Q(\rbzero.tex_r0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21214_ (.CLK(_00263_),
    .D(_01230_),
    .Q(\rbzero.tex_r0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21215_ (.CLK(_00264_),
    .D(_01231_),
    .Q(\rbzero.tex_r0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21216_ (.CLK(_00265_),
    .D(_01232_),
    .Q(\rbzero.tex_r0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21217_ (.CLK(_00266_),
    .D(_01233_),
    .Q(\rbzero.tex_r0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21218_ (.CLK(_00267_),
    .D(_01234_),
    .Q(\rbzero.tex_r0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21219_ (.CLK(_00268_),
    .D(_01235_),
    .Q(\rbzero.tex_r0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21220_ (.CLK(_00269_),
    .D(_01236_),
    .Q(\rbzero.tex_r0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21221_ (.CLK(_00270_),
    .D(_01237_),
    .Q(\rbzero.tex_r0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21222_ (.CLK(_00271_),
    .D(_01238_),
    .Q(\rbzero.tex_r0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21223_ (.CLK(_00272_),
    .D(_01239_),
    .Q(\rbzero.tex_r0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21224_ (.CLK(_00273_),
    .D(_01240_),
    .Q(\rbzero.tex_r1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21225_ (.CLK(_00274_),
    .D(_01241_),
    .Q(\rbzero.tex_r1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21226_ (.CLK(_00275_),
    .D(_01242_),
    .Q(\rbzero.tex_r1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21227_ (.CLK(_00276_),
    .D(_01243_),
    .Q(\rbzero.tex_r1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21228_ (.CLK(_00277_),
    .D(_01244_),
    .Q(\rbzero.tex_r1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21229_ (.CLK(_00278_),
    .D(_01245_),
    .Q(\rbzero.tex_r1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21230_ (.CLK(_00279_),
    .D(_01246_),
    .Q(\rbzero.tex_r1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21231_ (.CLK(_00280_),
    .D(_01247_),
    .Q(\rbzero.tex_r1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21232_ (.CLK(_00281_),
    .D(_01248_),
    .Q(\rbzero.tex_r1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21233_ (.CLK(_00282_),
    .D(_01249_),
    .Q(\rbzero.tex_r1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21234_ (.CLK(_00283_),
    .D(_01250_),
    .Q(\rbzero.tex_r1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21235_ (.CLK(_00284_),
    .D(_01251_),
    .Q(\rbzero.tex_r1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21236_ (.CLK(_00285_),
    .D(_01252_),
    .Q(\rbzero.tex_r1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21237_ (.CLK(_00286_),
    .D(_01253_),
    .Q(\rbzero.tex_r1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21238_ (.CLK(_00287_),
    .D(_01254_),
    .Q(\rbzero.tex_r1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21239_ (.CLK(_00288_),
    .D(_01255_),
    .Q(\rbzero.tex_r1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21240_ (.CLK(_00289_),
    .D(_01256_),
    .Q(\rbzero.tex_r1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21241_ (.CLK(_00290_),
    .D(_01257_),
    .Q(\rbzero.tex_r1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21242_ (.CLK(_00291_),
    .D(_01258_),
    .Q(\rbzero.tex_r1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21243_ (.CLK(_00292_),
    .D(_01259_),
    .Q(\rbzero.tex_r1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21244_ (.CLK(_00293_),
    .D(_01260_),
    .Q(\rbzero.tex_r1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21245_ (.CLK(_00294_),
    .D(_01261_),
    .Q(\rbzero.tex_r1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21246_ (.CLK(_00295_),
    .D(_01262_),
    .Q(\rbzero.tex_r1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21247_ (.CLK(_00296_),
    .D(_01263_),
    .Q(\rbzero.tex_r1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21248_ (.CLK(_00297_),
    .D(_01264_),
    .Q(\rbzero.tex_r1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21249_ (.CLK(_00298_),
    .D(_01265_),
    .Q(\rbzero.tex_r1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21250_ (.CLK(_00299_),
    .D(_01266_),
    .Q(\rbzero.tex_r1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21251_ (.CLK(_00300_),
    .D(_01267_),
    .Q(\rbzero.tex_r1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21252_ (.CLK(_00301_),
    .D(_01268_),
    .Q(\rbzero.tex_r1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21253_ (.CLK(_00302_),
    .D(_01269_),
    .Q(\rbzero.tex_r1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21254_ (.CLK(_00303_),
    .D(_01270_),
    .Q(\rbzero.tex_r1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21255_ (.CLK(_00304_),
    .D(_01271_),
    .Q(\rbzero.tex_r1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21256_ (.CLK(_00305_),
    .D(_01272_),
    .Q(\rbzero.tex_r1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21257_ (.CLK(_00306_),
    .D(_01273_),
    .Q(\rbzero.tex_r1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21258_ (.CLK(_00307_),
    .D(_01274_),
    .Q(\rbzero.tex_r1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21259_ (.CLK(_00308_),
    .D(_01275_),
    .Q(\rbzero.tex_r1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21260_ (.CLK(_00309_),
    .D(_01276_),
    .Q(\rbzero.tex_r1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21261_ (.CLK(_00310_),
    .D(_01277_),
    .Q(\rbzero.tex_r1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21262_ (.CLK(_00311_),
    .D(_01278_),
    .Q(\rbzero.tex_r1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21263_ (.CLK(_00312_),
    .D(_01279_),
    .Q(\rbzero.tex_r1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21264_ (.CLK(_00313_),
    .D(_01280_),
    .Q(\rbzero.tex_r1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21265_ (.CLK(_00314_),
    .D(_01281_),
    .Q(\rbzero.tex_r1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21266_ (.CLK(_00315_),
    .D(_01282_),
    .Q(\rbzero.tex_r1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21267_ (.CLK(_00316_),
    .D(_01283_),
    .Q(\rbzero.tex_r1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21268_ (.CLK(_00317_),
    .D(_01284_),
    .Q(\rbzero.tex_r1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21269_ (.CLK(_00318_),
    .D(_01285_),
    .Q(\rbzero.tex_r1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21270_ (.CLK(_00319_),
    .D(_01286_),
    .Q(\rbzero.tex_r1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21271_ (.CLK(_00320_),
    .D(_01287_),
    .Q(\rbzero.tex_r1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21272_ (.CLK(_00321_),
    .D(_01288_),
    .Q(\rbzero.tex_r1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21273_ (.CLK(_00322_),
    .D(_01289_),
    .Q(\rbzero.tex_r1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21274_ (.CLK(_00323_),
    .D(_01290_),
    .Q(\rbzero.tex_r1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21275_ (.CLK(_00324_),
    .D(_01291_),
    .Q(\rbzero.tex_r1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21276_ (.CLK(_00325_),
    .D(_01292_),
    .Q(\rbzero.tex_r1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21277_ (.CLK(_00326_),
    .D(_01293_),
    .Q(\rbzero.tex_r1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21278_ (.CLK(_00327_),
    .D(_01294_),
    .Q(\rbzero.tex_r1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21279_ (.CLK(_00328_),
    .D(_01295_),
    .Q(\rbzero.tex_r1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21280_ (.CLK(_00329_),
    .D(_01296_),
    .Q(\rbzero.tex_r1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21281_ (.CLK(_00330_),
    .D(_01297_),
    .Q(\rbzero.tex_r1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21282_ (.CLK(_00331_),
    .D(_01298_),
    .Q(\rbzero.tex_r1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21283_ (.CLK(_00332_),
    .D(_01299_),
    .Q(\rbzero.tex_r1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21284_ (.CLK(_00333_),
    .D(_01300_),
    .Q(\rbzero.tex_r1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21285_ (.CLK(_00334_),
    .D(_01301_),
    .Q(\rbzero.tex_r1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21286_ (.CLK(_00335_),
    .D(_01302_),
    .Q(\rbzero.tex_r1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21287_ (.CLK(_00336_),
    .D(_01303_),
    .Q(\rbzero.tex_r1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21288_ (.CLK(net114),
    .D(_01304_),
    .Q(\gpout5.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21289_ (.CLK(net114),
    .D(_01305_),
    .Q(\gpout5.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21290_ (.CLK(net133),
    .D(_01306_),
    .Q(\rbzero.texV[-12] ));
 sky130_fd_sc_hd__dfxtp_1 _21291_ (.CLK(net134),
    .D(_01307_),
    .Q(\rbzero.texV[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21292_ (.CLK(net134),
    .D(_01308_),
    .Q(\rbzero.texV[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21293_ (.CLK(net134),
    .D(_01309_),
    .Q(\rbzero.texV[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21294_ (.CLK(net134),
    .D(_01310_),
    .Q(\rbzero.texV[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21295_ (.CLK(net134),
    .D(_01311_),
    .Q(\rbzero.texV[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21296_ (.CLK(net134),
    .D(_01312_),
    .Q(\rbzero.texV[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21297_ (.CLK(net134),
    .D(_01313_),
    .Q(\rbzero.texV[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21298_ (.CLK(net114),
    .D(_01314_),
    .Q(\rbzero.texV[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21299_ (.CLK(net133),
    .D(_01315_),
    .Q(\rbzero.texV[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21300_ (.CLK(net134),
    .D(_01316_),
    .Q(\rbzero.texV[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21301_ (.CLK(net132),
    .D(_01317_),
    .Q(\rbzero.texV[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21302_ (.CLK(net128),
    .D(_01318_),
    .Q(\rbzero.texV[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21303_ (.CLK(net127),
    .D(_01319_),
    .Q(\rbzero.texV[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21304_ (.CLK(net128),
    .D(_01320_),
    .Q(\rbzero.texV[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21305_ (.CLK(net129),
    .D(_01321_),
    .Q(\rbzero.texV[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21306_ (.CLK(net132),
    .D(_01322_),
    .Q(\rbzero.texV[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21307_ (.CLK(net133),
    .D(_01323_),
    .Q(\rbzero.texV[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21308_ (.CLK(net114),
    .D(_01324_),
    .Q(\rbzero.texV[6] ));
 sky130_fd_sc_hd__dfxtp_2 _21309_ (.CLK(net114),
    .D(_01325_),
    .Q(\rbzero.texV[7] ));
 sky130_fd_sc_hd__dfxtp_2 _21310_ (.CLK(net112),
    .D(_01326_),
    .Q(\rbzero.texV[8] ));
 sky130_fd_sc_hd__dfxtp_2 _21311_ (.CLK(net112),
    .D(_01327_),
    .Q(\rbzero.texV[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21312_ (.CLK(net111),
    .D(_01328_),
    .Q(\rbzero.texV[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21313_ (.CLK(net111),
    .D(_01329_),
    .Q(\rbzero.texV[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21314_ (.CLK(_00337_),
    .D(_01330_),
    .Q(\rbzero.tex_b1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21315_ (.CLK(_00338_),
    .D(_01331_),
    .Q(\rbzero.tex_b1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21316_ (.CLK(_00339_),
    .D(_01332_),
    .Q(\rbzero.tex_b1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21317_ (.CLK(_00340_),
    .D(_01333_),
    .Q(\rbzero.tex_b1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21318_ (.CLK(_00341_),
    .D(_01334_),
    .Q(\rbzero.tex_b1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21319_ (.CLK(_00342_),
    .D(_01335_),
    .Q(\rbzero.tex_b1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21320_ (.CLK(_00343_),
    .D(_01336_),
    .Q(\rbzero.tex_b1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21321_ (.CLK(_00344_),
    .D(_01337_),
    .Q(\rbzero.tex_b1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21322_ (.CLK(_00345_),
    .D(_01338_),
    .Q(\rbzero.tex_b1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21323_ (.CLK(_00346_),
    .D(_01339_),
    .Q(\rbzero.tex_b1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21324_ (.CLK(_00347_),
    .D(_01340_),
    .Q(\rbzero.tex_b1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21325_ (.CLK(_00348_),
    .D(_01341_),
    .Q(\rbzero.tex_b1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21326_ (.CLK(_00349_),
    .D(_01342_),
    .Q(\rbzero.tex_b1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21327_ (.CLK(_00350_),
    .D(_01343_),
    .Q(\rbzero.tex_b1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21328_ (.CLK(_00351_),
    .D(_01344_),
    .Q(\rbzero.tex_b1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21329_ (.CLK(_00352_),
    .D(_01345_),
    .Q(\rbzero.tex_b1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21330_ (.CLK(_00353_),
    .D(_01346_),
    .Q(\rbzero.tex_b1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21331_ (.CLK(_00354_),
    .D(_01347_),
    .Q(\rbzero.tex_b1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21332_ (.CLK(_00355_),
    .D(_01348_),
    .Q(\rbzero.tex_b1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21333_ (.CLK(_00356_),
    .D(_01349_),
    .Q(\rbzero.tex_b1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21334_ (.CLK(_00357_),
    .D(_01350_),
    .Q(\rbzero.tex_b1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21335_ (.CLK(_00358_),
    .D(_01351_),
    .Q(\rbzero.tex_b1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21336_ (.CLK(_00359_),
    .D(_01352_),
    .Q(\rbzero.tex_b1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21337_ (.CLK(_00360_),
    .D(_01353_),
    .Q(\rbzero.tex_b1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21338_ (.CLK(_00361_),
    .D(_01354_),
    .Q(\rbzero.tex_b1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21339_ (.CLK(_00362_),
    .D(_01355_),
    .Q(\rbzero.tex_b1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21340_ (.CLK(_00363_),
    .D(_01356_),
    .Q(\rbzero.tex_b1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21341_ (.CLK(_00364_),
    .D(_01357_),
    .Q(\rbzero.tex_b1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21342_ (.CLK(_00365_),
    .D(_01358_),
    .Q(\rbzero.tex_b1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21343_ (.CLK(_00366_),
    .D(_01359_),
    .Q(\rbzero.tex_b1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21344_ (.CLK(_00367_),
    .D(_01360_),
    .Q(\rbzero.tex_b1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21345_ (.CLK(_00368_),
    .D(_01361_),
    .Q(\rbzero.tex_b1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21346_ (.CLK(_00369_),
    .D(_01362_),
    .Q(\rbzero.tex_b1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21347_ (.CLK(_00370_),
    .D(_01363_),
    .Q(\rbzero.tex_b1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21348_ (.CLK(_00371_),
    .D(_01364_),
    .Q(\rbzero.tex_b1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21349_ (.CLK(_00372_),
    .D(_01365_),
    .Q(\rbzero.tex_b1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21350_ (.CLK(_00373_),
    .D(_01366_),
    .Q(\rbzero.tex_b1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21351_ (.CLK(_00374_),
    .D(_01367_),
    .Q(\rbzero.tex_b1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21352_ (.CLK(_00375_),
    .D(_01368_),
    .Q(\rbzero.tex_b1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21353_ (.CLK(_00376_),
    .D(_01369_),
    .Q(\rbzero.tex_b1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21354_ (.CLK(_00377_),
    .D(_01370_),
    .Q(\rbzero.tex_b1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21355_ (.CLK(_00378_),
    .D(_01371_),
    .Q(\rbzero.tex_b1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21356_ (.CLK(_00379_),
    .D(_01372_),
    .Q(\rbzero.tex_b1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21357_ (.CLK(_00380_),
    .D(_01373_),
    .Q(\rbzero.tex_b1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21358_ (.CLK(_00381_),
    .D(_01374_),
    .Q(\rbzero.tex_b1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21359_ (.CLK(_00382_),
    .D(_01375_),
    .Q(\rbzero.tex_b1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21360_ (.CLK(_00383_),
    .D(_01376_),
    .Q(\rbzero.tex_b1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21361_ (.CLK(_00384_),
    .D(_01377_),
    .Q(\rbzero.tex_b1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21362_ (.CLK(_00385_),
    .D(_01378_),
    .Q(\rbzero.tex_b1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21363_ (.CLK(_00386_),
    .D(_01379_),
    .Q(\rbzero.tex_b1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21364_ (.CLK(_00387_),
    .D(_01380_),
    .Q(\rbzero.tex_b1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21365_ (.CLK(_00388_),
    .D(_01381_),
    .Q(\rbzero.tex_b1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21366_ (.CLK(_00389_),
    .D(_01382_),
    .Q(\rbzero.tex_b1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21367_ (.CLK(_00390_),
    .D(_01383_),
    .Q(\rbzero.tex_b1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21368_ (.CLK(_00391_),
    .D(_01384_),
    .Q(\rbzero.tex_b1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21369_ (.CLK(_00392_),
    .D(_01385_),
    .Q(\rbzero.tex_b1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21370_ (.CLK(_00393_),
    .D(_01386_),
    .Q(\rbzero.tex_b1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21371_ (.CLK(_00394_),
    .D(_01387_),
    .Q(\rbzero.tex_b1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21372_ (.CLK(_00395_),
    .D(_01388_),
    .Q(\rbzero.tex_b1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21373_ (.CLK(_00396_),
    .D(_01389_),
    .Q(\rbzero.tex_b1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21374_ (.CLK(_00397_),
    .D(_01390_),
    .Q(\rbzero.tex_b1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21375_ (.CLK(_00398_),
    .D(_01391_),
    .Q(\rbzero.tex_b1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21376_ (.CLK(_00399_),
    .D(_01392_),
    .Q(\rbzero.tex_b1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21377_ (.CLK(_00400_),
    .D(_01393_),
    .Q(\rbzero.tex_b1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21378_ (.CLK(net119),
    .D(_01394_),
    .Q(\rbzero.traced_texVinit[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21379_ (.CLK(net127),
    .D(_01395_),
    .Q(\rbzero.traced_texVinit[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21380_ (.CLK(net127),
    .D(_01396_),
    .Q(\rbzero.traced_texVinit[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21381_ (.CLK(net97),
    .D(_01397_),
    .Q(\rbzero.traced_texVinit[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21382_ (.CLK(net113),
    .D(_01398_),
    .Q(\rbzero.traced_texVinit[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21383_ (.CLK(net112),
    .D(_01399_),
    .Q(\rbzero.traced_texVinit[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21384_ (.CLK(net112),
    .D(_01400_),
    .Q(\rbzero.traced_texVinit[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21385_ (.CLK(net113),
    .D(_01401_),
    .Q(\rbzero.traced_texVinit[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21386_ (.CLK(net109),
    .D(_01402_),
    .Q(\rbzero.traced_texVinit[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21387_ (.CLK(net109),
    .D(_01403_),
    .Q(\rbzero.traced_texVinit[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21388_ (.CLK(net109),
    .D(_01404_),
    .Q(\rbzero.traced_texVinit[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21389_ (.CLK(net109),
    .D(_01405_),
    .Q(\rbzero.traced_texVinit[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21390_ (.CLK(net110),
    .D(_01406_),
    .Q(\gpout0.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21391_ (.CLK(net110),
    .D(_01407_),
    .Q(\gpout0.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21392_ (.CLK(net114),
    .D(_01408_),
    .Q(\gpout1.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21393_ (.CLK(net108),
    .D(_01409_),
    .Q(\gpout1.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21394_ (.CLK(net86),
    .D(_01410_),
    .Q(\rbzero.wall_tracer.rayAddendX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21395_ (.CLK(net86),
    .D(_01411_),
    .Q(\rbzero.wall_tracer.rayAddendX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21396_ (.CLK(net86),
    .D(_01412_),
    .Q(\rbzero.wall_tracer.rayAddendX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21397_ (.CLK(net86),
    .D(_01413_),
    .Q(\rbzero.wall_tracer.rayAddendX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21398_ (.CLK(net83),
    .D(_01414_),
    .Q(\rbzero.wall_tracer.rayAddendY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21399_ (.CLK(net83),
    .D(_01415_),
    .Q(\rbzero.wall_tracer.rayAddendY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21400_ (.CLK(net86),
    .D(_01416_),
    .Q(\rbzero.wall_tracer.rayAddendY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21401_ (.CLK(net86),
    .D(_01417_),
    .Q(\rbzero.wall_tracer.rayAddendY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21402_ (.CLK(net110),
    .D(_01418_),
    .Q(\gpout2.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21403_ (.CLK(net106),
    .D(_01419_),
    .Q(\gpout2.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21404_ (.CLK(net114),
    .D(_01420_),
    .Q(\gpout3.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21405_ (.CLK(net114),
    .D(_01421_),
    .Q(\gpout3.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21406_ (.CLK(net115),
    .D(_01422_),
    .Q(\gpout4.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21407_ (.CLK(net115),
    .D(_01423_),
    .Q(\gpout4.clk_div[1] ));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_143 (.LO(net143));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_144 (.LO(net144));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_145 (.LO(net145));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_146 (.LO(net146));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_147 (.LO(net147));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_148 (.LO(net148));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_149 (.LO(net149));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_150 (.LO(net150));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_151 (.LO(net151));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_152 (.LO(net152));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_153 (.LO(net153));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_154 (.LO(net154));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_155 (.LO(net155));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_156 (.LO(net156));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_157 (.LO(net157));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_158 (.LO(net158));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_159 (.LO(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_01823_));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__buf_6 input1 (.A(i_clk),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input2 (.A(i_debug_vec_overlay),
    .X(net2));
 sky130_fd_sc_hd__buf_6 input3 (.A(i_gpout0_sel[0]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(i_gpout0_sel[1]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(i_gpout0_sel[2]),
    .X(net5));
 sky130_fd_sc_hd__buf_6 input6 (.A(i_gpout0_sel[3]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(i_gpout0_sel[4]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(i_gpout0_sel[5]),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input9 (.A(i_gpout1_sel[0]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 input10 (.A(i_gpout1_sel[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(i_gpout1_sel[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(i_gpout1_sel[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_8 input13 (.A(i_gpout1_sel[4]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(i_gpout1_sel[5]),
    .X(net14));
 sky130_fd_sc_hd__buf_6 input15 (.A(i_gpout2_sel[0]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_8 input16 (.A(i_gpout2_sel[1]),
    .X(net16));
 sky130_fd_sc_hd__buf_6 input17 (.A(i_gpout2_sel[2]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input18 (.A(i_gpout2_sel[3]),
    .X(net18));
 sky130_fd_sc_hd__buf_6 input19 (.A(i_gpout2_sel[4]),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input20 (.A(i_gpout2_sel[5]),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input21 (.A(i_gpout3_sel[0]),
    .X(net21));
 sky130_fd_sc_hd__buf_4 input22 (.A(i_gpout3_sel[1]),
    .X(net22));
 sky130_fd_sc_hd__buf_4 input23 (.A(i_gpout3_sel[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_8 input24 (.A(i_gpout3_sel[3]),
    .X(net24));
 sky130_fd_sc_hd__buf_4 input25 (.A(i_gpout3_sel[4]),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(i_gpout3_sel[5]),
    .X(net26));
 sky130_fd_sc_hd__buf_6 input27 (.A(i_gpout4_sel[0]),
    .X(net27));
 sky130_fd_sc_hd__buf_6 input28 (.A(i_gpout4_sel[1]),
    .X(net28));
 sky130_fd_sc_hd__buf_4 input29 (.A(i_gpout4_sel[2]),
    .X(net29));
 sky130_fd_sc_hd__buf_6 input30 (.A(i_gpout4_sel[3]),
    .X(net30));
 sky130_fd_sc_hd__buf_4 input31 (.A(i_gpout4_sel[4]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(i_gpout4_sel[5]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 input33 (.A(i_gpout5_sel[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(i_gpout5_sel[1]),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(i_gpout5_sel[2]),
    .X(net35));
 sky130_fd_sc_hd__buf_4 input36 (.A(i_gpout5_sel[3]),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(i_gpout5_sel[4]),
    .X(net37));
 sky130_fd_sc_hd__buf_6 input38 (.A(i_gpout5_sel[5]),
    .X(net38));
 sky130_fd_sc_hd__buf_6 input39 (.A(i_mode[0]),
    .X(net39));
 sky130_fd_sc_hd__buf_8 input40 (.A(i_mode[1]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_8 input41 (.A(i_mode[2]),
    .X(net41));
 sky130_fd_sc_hd__buf_8 input42 (.A(i_reg_csb),
    .X(net42));
 sky130_fd_sc_hd__buf_6 input43 (.A(i_reg_mosi),
    .X(net43));
 sky130_fd_sc_hd__buf_6 input44 (.A(i_reg_sclk),
    .X(net44));
 sky130_fd_sc_hd__buf_8 input45 (.A(i_reset_lock_a),
    .X(net45));
 sky130_fd_sc_hd__buf_8 input46 (.A(i_reset_lock_b),
    .X(net46));
 sky130_fd_sc_hd__buf_6 input47 (.A(i_tex_in[0]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(i_tex_in[1]),
    .X(net48));
 sky130_fd_sc_hd__buf_4 input49 (.A(i_tex_in[2]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 input50 (.A(i_tex_in[3]),
    .X(net50));
 sky130_fd_sc_hd__buf_4 input51 (.A(i_vec_csb),
    .X(net51));
 sky130_fd_sc_hd__buf_8 input52 (.A(i_vec_mosi),
    .X(net52));
 sky130_fd_sc_hd__buf_6 input53 (.A(i_vec_sclk),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 fanout54 (.A(net59),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 fanout55 (.A(net57),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 fanout56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 fanout57 (.A(net58),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 fanout58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout59 (.A(net73),
    .X(net59));
 sky130_fd_sc_hd__buf_2 fanout60 (.A(net73),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 fanout61 (.A(net73),
    .X(net61));
 sky130_fd_sc_hd__buf_2 fanout62 (.A(net64),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 fanout63 (.A(net64),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout64 (.A(net72),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 fanout65 (.A(net72),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 fanout66 (.A(net72),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 fanout67 (.A(net69),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 fanout68 (.A(net69),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 fanout69 (.A(net72),
    .X(net69));
 sky130_fd_sc_hd__buf_2 fanout70 (.A(net72),
    .X(net70));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout71 (.A(net72),
    .X(net71));
 sky130_fd_sc_hd__buf_2 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_4 fanout73 (.A(net1),
    .X(net73));
 sky130_fd_sc_hd__buf_2 fanout74 (.A(net77),
    .X(net74));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout75 (.A(net77),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 fanout76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 fanout77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout78 (.A(net1),
    .X(net78));
 sky130_fd_sc_hd__buf_2 fanout79 (.A(net80),
    .X(net79));
 sky130_fd_sc_hd__buf_2 fanout80 (.A(net83),
    .X(net80));
 sky130_fd_sc_hd__buf_2 fanout81 (.A(net83),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 fanout82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 fanout83 (.A(net98),
    .X(net83));
 sky130_fd_sc_hd__buf_2 fanout84 (.A(net89),
    .X(net84));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__buf_2 fanout86 (.A(net89),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 fanout87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 fanout88 (.A(net89),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 fanout89 (.A(net98),
    .X(net89));
 sky130_fd_sc_hd__buf_2 fanout90 (.A(net92),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 fanout91 (.A(net92),
    .X(net91));
 sky130_fd_sc_hd__buf_2 fanout92 (.A(net98),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__buf_2 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__buf_2 fanout95 (.A(net98),
    .X(net95));
 sky130_fd_sc_hd__buf_2 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 fanout97 (.A(net98),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 fanout98 (.A(net141),
    .X(net98));
 sky130_fd_sc_hd__buf_2 fanout99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__buf_2 fanout100 (.A(net104),
    .X(net100));
 sky130_fd_sc_hd__buf_2 fanout101 (.A(net104),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 fanout102 (.A(net104),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 fanout103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__buf_2 fanout104 (.A(net108),
    .X(net104));
 sky130_fd_sc_hd__buf_2 fanout105 (.A(net108),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 fanout106 (.A(net108),
    .X(net106));
 sky130_fd_sc_hd__buf_2 fanout107 (.A(net108),
    .X(net107));
 sky130_fd_sc_hd__buf_2 fanout108 (.A(net141),
    .X(net108));
 sky130_fd_sc_hd__buf_2 fanout109 (.A(net115),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 fanout110 (.A(net115),
    .X(net110));
 sky130_fd_sc_hd__buf_2 fanout111 (.A(net113),
    .X(net111));
 sky130_fd_sc_hd__buf_2 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 fanout113 (.A(net115),
    .X(net113));
 sky130_fd_sc_hd__buf_2 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 fanout115 (.A(net141),
    .X(net115));
 sky130_fd_sc_hd__buf_2 fanout116 (.A(net122),
    .X(net116));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout117 (.A(net122),
    .X(net117));
 sky130_fd_sc_hd__buf_2 fanout118 (.A(net122),
    .X(net118));
 sky130_fd_sc_hd__buf_2 fanout119 (.A(net122),
    .X(net119));
 sky130_fd_sc_hd__buf_2 fanout120 (.A(net122),
    .X(net120));
 sky130_fd_sc_hd__buf_2 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__buf_2 fanout122 (.A(net126),
    .X(net122));
 sky130_fd_sc_hd__buf_2 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 fanout126 (.A(net141),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 fanout127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__buf_2 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 fanout129 (.A(net140),
    .X(net129));
 sky130_fd_sc_hd__buf_2 fanout130 (.A(net140),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 fanout131 (.A(net140),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 fanout132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__buf_2 fanout134 (.A(net140),
    .X(net134));
 sky130_fd_sc_hd__buf_2 fanout135 (.A(net139),
    .X(net135));
 sky130_fd_sc_hd__buf_2 fanout136 (.A(net139),
    .X(net136));
 sky130_fd_sc_hd__buf_2 fanout137 (.A(net139),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_2 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__buf_2 fanout140 (.A(net141),
    .X(net140));
 sky130_fd_sc_hd__buf_4 fanout141 (.A(net1),
    .X(net141));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_142 (.LO(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_01823_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_02720_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_07189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_09200_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_09470_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(o_rgb[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(o_rgb[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(o_rgb[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\rbzero.pov.mosi ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\rbzero.traced_texa[-11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\rbzero.wall_tracer.visualWallDist[-3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\rbzero.wall_tracer.visualWallDist[-5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_07172_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_07838_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_10056_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(o_rgb[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\rbzero.wall_tracer.visualWallDist[-9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\rbzero.wall_tracer.visualWallDist[-9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_02708_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1092 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1487 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1176 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1250 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1246 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1234 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1247 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1223 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1274 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1274 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1265 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1271 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1319 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1280 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1274 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1176 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1299 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1207 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1224 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1278 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1262 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_919 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1204 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_843 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1143 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_919 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1207 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1178 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1226 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1178 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_843 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1191 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1120 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1208 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1246 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1180 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1246 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1250 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1066 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1278 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1250 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1242 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1208 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1222 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1234 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1242 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1148 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1066 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_1492 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_1490 ();
 assign o_rgb[0] = net142;
 assign o_rgb[10] = net150;
 assign o_rgb[11] = net151;
 assign o_rgb[12] = net152;
 assign o_rgb[13] = net153;
 assign o_rgb[16] = net154;
 assign o_rgb[17] = net155;
 assign o_rgb[18] = net156;
 assign o_rgb[19] = net157;
 assign o_rgb[1] = net143;
 assign o_rgb[20] = net158;
 assign o_rgb[21] = net159;
 assign o_rgb[2] = net144;
 assign o_rgb[3] = net145;
 assign o_rgb[4] = net146;
 assign o_rgb[5] = net147;
 assign o_rgb[8] = net148;
 assign o_rgb[9] = net149;
endmodule

